// THIS FILE IS WRITTEN IN SJIS CODE SET

import_C( "tecs.h" );

// '�\' �̑��o�C�g�� 0x5c (�o�b�N�X���b�V�� '\')�ŁA'"' �̒��O�ɂ���ƁA
// �����񃊃e���������Ă��Ȃ����̂悤�Ɍ�F�����\��������

const char_t * const PtrConst = "�~�\";

signature sSig {
	ER  func( [in]int32_t par );
};

celltype tCelltype {
	attr {
		char_t *StrPtr = "�w�\";
		int32_t a = '�\';
		int32_t b = '��';
		int32_t c = '\n';
	};
	entry sSig eEnt;

	factory {
		write( "tecsgen.cfg", "�~�\%s", StrPtr );
	};
};

cell tCelltype Cell {
};
