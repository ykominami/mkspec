/*
 *                        +------------------------------------------------------------------+
 *                        |   +---------------------------+   +---------------------------+  |
 *  +-----------------+   |   |   +--------+  +--------+  | s3|   +--------+  +--------+  |  |  +-------------+
 *  |                 | s1|   |   |        |s2|        |--+---|>--|>       |s4|        |  |  |s5|             |
 *  |  Cell_clnt c[0] |-+-|---|>--|> Cell1 |--|> Cell2 |  | sB|   | Cell3  |--|> Cell4 |--+--|--|> Cell_serv1 |
 *  |            c[1] |-+ |   |   |        |  |       <|-<|---+---|        |  |        |  |  |  |             |
 *  +-----------------+ | |   |   +--------+  +--------+  |   |   +--------+  +--------+  |  |  +-------------+
 *                      | |   |       tComp11 comp11      |   |       tComp12 comp12      |  |
 *                      | |   +---------------------------+   +---------------------------+  |
 *                      | |                          tComp3 Comp1                            |
 *                      | +------------------------------------------------------------------+
 *                      |
 *                      | +------------------------------------------------------------------+
 *                      | |   +---------------------------+   +---------------------------+  |
 *                      | |   |   +--------+  +--------+  | s3|   +--------+  +--------+  |  |  +-------------+
 *                      | |   |   |        |s2|        |--+---|>--|>       |s4|        |  |  |s5|             |
 *                      +-|>--|>--|> Cell1 |--|> Cell2 |  | sB|   |  Cell3 |--|> Cell4 |--+--|--|> Cell_serv2 |
 *                        |   |   |        |  |       <|-<|---+---|        |  |        |  |  |  |             |
 *                        |   |   +--------+  +--------+  |   |   +--------+  +--------+  |  |  +-------------+
 *                        |   |       tComp11 comp11      |   |       tComp12 comp12      |  |
 *                        |   +---------------------------+   +---------------------------+  |
 *                        |                          tComp3 Comp2                            |
 *                        +------------------------------------------------------------------+
 */
import_C( "tecs.h" );
import( <cygwin_kernel.cdl> );

signature sSig1 {
  int32_t  func1( [in]int32_t a );
  int32_t  func2( [in]int32_t a );
};

signature sSig2 {
  int32_t  func1( [in]int32_t a );
  int32_t  func2( [in]int32_t a );
};

signature sSig3 {
  int32_t  func1( [in]int32_t a );
  int32_t  func2( [in]int32_t a );
};

signature sSig4 {
  int32_t  func1( [in]int32_t a );
  int32_t  func2( [in]int32_t a );
};

signature sSig5 {
  int32_t  func1( [in]int32_t a );
  int32_t  func2( [in]int32_t a );
};

signature sSigB {
  int32_t  func1( [in]int32_t a );
  int32_t  func2( [in]int32_t a );
};


celltype tCell1 {
    entry sSig1 eEntry1;
    call  sSig2 cCall1;
    attr{
        char *name = C_EXP( "\"$cell$\"" );
        int32_t a;
    };
};

celltype tCell2 {
    entry sSig2 eEntry2;
    call  sSig3 cCall2[2];
    entry sSigB eEntryB;
    attr{
        char *name = C_EXP( "\"$cell$\"" );
        int32_t a;
    };
};

composite tComp11 {
    call sSig3 cCall[2];
    entry sSig1 eEntry;
    entry sSigB eEntryB;

    cell tCell1 cell1{
        cCall1 = cell2.eEntry2;
        a = 10;
    };
    cell tCell2 cell2 {
        cCall2 => cCall;
        a = 20;
    };

    eEntry  => cell1.eEntry1;
    eEntryB => cell2.eEntryB;
};


celltype tCell3 {
    entry sSig3 eEntry3[2];
    call  sSig4 cCall3;
    call  sSigB cCallB;
    attr{
        char *name = C_EXP( "\"$cell$\"" );
        int32_t a;
    };
};

celltype tCell4 {
    entry sSig4 eEntry4;
    call  sSig5 cCall4;
    attr{
        char *name = C_EXP( "\"$cell$\"" );
        int32_t a;
    };
};

composite tComp12 {

  attr {
    int32_t a = 40;
  };
  call sSig5 cCall;
  call sSigB cCallB;
  entry sSig3 eEntry[2];

  cell tCell4 cell4;

  cell tCell3 cell3{
    cCall3 = cell4.eEntry4;
    cCallB => composite.cCallB;
    a = 30;
  };
  cell tCell4 cell4 {
    cCall4 => cCall;
    a = composite.a;
  };

  eEntry => cell3.eEntry3;
};


composite tComp3 {

  attr {
    int32_t a;
  };
  call sSig5 cCall;
  entry sSig1 eEntry;

  cell tComp12 comp12;

  cell tComp11 comp11 {
    cCall[] = comp12.eEntry[1];
    cCall[] = comp12.eEntry[0];
  };

  cell tComp12 comp12 {
    cCallB = comp11.eEntryB;
    cCall => composite.cCall;
    a = composite.a;
  };

  eEntry => comp11.eEntry;
};

celltype tCell_serv {
  entry sSig5 eEntry;
  attr {
    int32_t a;
  };
};

celltype tCell_clnt {
  entry sTaskBody eMain;
  call sSig1 cCall[];
  attr {
    int32_t a;
  };
};

cell tTask Task1 {
  cTaskBody = cell_clnt.eMain;
  priority = 0;
  stackSize = 4096;
  attribute = C_EXP( "TA_ACT" );
//  attribute = C_EXP( "TA_NULL" );
};
cell tCell_clnt cell_clnt {
  a = 30;
  cCall[0] = comp1.eEntry;
  cCall[1] = comp2.eEntry;
  cCall[2] = rLargeComp::LargeComp.eServ1;
  cCall[3] = rLargeComp::LargeComp.eServ2;
};

cell tComp3 comp2 {
  a=10;
  cCall = cell_serv2.eEntry;
};

cell tCell_serv cell_serv2{
   a = 201;
};

cell tComp3 comp1 {
  a=101;
  cCall = cell_serv1.eEntry;
};

cell tCell_serv cell_serv1{
   a = 5;
};

//////////    ///////////
composite tLargeComp {
  entry  sSig1  eServ1;
  entry  sSig1  eServ2;
  call   sSig5 cCall1;
  call   sSig5 cCall2;

  cell tComp3 comp1 {
    a=101;
    cCall => composite.cCall1;
  };
  cell tComp3 comp2 {
    a=10;
    cCall => composite.cCall2;
  };
  composite.eServ1 => comp1.eEntry;
  composite.eServ2 => comp2.eEntry;
};

[in_through()]
region rLargeComp {
/*  cell tTask Task2{
    cBody = CellClnt.eMain;
    priority = 0;
    stackSize = 4096;
//    attribute = C_EXP( "TA_NULL" );
    attribute = C_EXP( "TA_ACT" );
  };

  cell tCell_clnt CellClnt{
    cCall[0] = LargeComp.eServ1;
    cCall[1] = LargeComp.eServ2;
    a = 102;
  };
*/
  cell tLargeComp LargeComp {
    cCall1 = CellServ1.eEntry;
    cCall2 = CellServ2.eEntry;
  };

  cell tCell_serv CellServ1{
    a = 5;
  };
  
  cell tCell_serv CellServ2{
    a = 201;
  };
};

