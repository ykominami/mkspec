/*------------ TECSInfoPlugin post code ------------*/
region rTEMP{
    region rTECSInfo {

        /*** :: namespace information cell ***/
        cell nTECSInfo::tNamespaceInfo _RootNamespaceInfo{
            name = "::";

            /* SIGNATURE info */
            cSignatureInfo[] = sTaskBodySignatureInfo.eSignatureInfo;
            cSignatureInfo[] = sTaskExceptionBodySignatureInfo.eSignatureInfo;
            cSignatureInfo[] = sTaskSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = sKernelSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = siKernelSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = sSemaphoreSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = siSemaphoreSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = sEventflagSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = siEventflagSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = sDataqueueSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = siDataqueueSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = sPutStringSignatureInfo.eSignatureInfo;

            /* CELLTYPE info */
            cCelltypeInfo[] = tTaskCelltypeInfo.eCelltypeInfo;
            cCelltypeInfo[] = tPutStringStdioCelltypeInfo.eCelltypeInfo;
            cCelltypeInfo[] = tHelloWorldCelltypeInfo.eCelltypeInfo;
            cCelltypeInfo[] = tTaskMainCelltypeInfo.eCelltypeInfo;

            /* NAMESPACE info */
            cNamespaceInfo[] = nTECSInfoNamespaceInfo.eNamespaceInfo;
        };   /* cell nTECSInfo::tNamespaceInfo _RootNamespaceInfo */

        /*** sTaskBody signature information ****/
        cell nTECSInfo::tSignatureInfo sTaskBodySignatureInfo {
            name            = "sTaskBody";
            cFunctionInfo[] = sTaskBody_mainFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo sTaskBody_mainFunctionInfo {
            name            = "main";
            bOneway         = false;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };

        /*** sTaskExceptionBody signature information ****/
        cell nTECSInfo::tSignatureInfo sTaskExceptionBodySignatureInfo {
            name            = "sTaskExceptionBody";
            cFunctionInfo[] = sTaskExceptionBody_mainFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo sTaskExceptionBody_mainFunctionInfo {
            name            = "main";
            bOneway         = false;
            cParamInfo[]    = sTaskExceptionBody_main_patternParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sTaskExceptionBody_main_patternParamInfo {
            name            = "pattern";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = TEXPTNTypeInfo.eTypeInfo;
        };

        /*** sTask signature information ****/
        cell nTECSInfo::tSignatureInfo sTaskSignatureInfo {
            name            = "sTask";
            cFunctionInfo[] = sTask_activateFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sTask_suspendFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sTask_resumeFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo sTask_activateFunctionInfo {
            name            = "activate";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sTask_suspendFunctionInfo {
            name            = "suspend";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sTask_resumeFunctionInfo {
            name            = "resume";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };

        /*** sKernel signature information ****/
        cell nTECSInfo::tSignatureInfo sKernelSignatureInfo {
            name            = "sKernel";
            cFunctionInfo[] = sKernel_delayFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sKernel_exitTaskFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sKernel_getTimeFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sKernel_getMicroTimeFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sKernel_exitKernelFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo sKernel_delayFunctionInfo {
            name            = "delay";
            bOneway         = false;
            cParamInfo[]    = sKernel_delay_delay_timeParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sKernel_delay_delay_timeParamInfo {
            name            = "delay_time";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = RELTIMTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sKernel_exitTaskFunctionInfo {
            name            = "exitTask";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sKernel_getTimeFunctionInfo {
            name            = "getTime";
            bOneway         = false;
            cParamInfo[]    = sKernel_getTime_p_system_timeParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sKernel_getTime_p_system_timeParamInfo {
            name            = "p_system_time";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = SYSTIM_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sKernel_getMicroTimeFunctionInfo {
            name            = "getMicroTime";
            bOneway         = false;
            cParamInfo[]    = sKernel_getMicroTime_p_system_micro_timeParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sKernel_getMicroTime_p_system_micro_timeParamInfo {
            name            = "p_system_micro_time";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = SYSUTM_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sKernel_exitKernelFunctionInfo {
            name            = "exitKernel";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };

        /*** siKernel signature information ****/
        cell nTECSInfo::tSignatureInfo siKernelSignatureInfo {
            name            = "siKernel";
            cFunctionInfo[] = siKernel_getMicroTimeFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo siKernel_getMicroTimeFunctionInfo {
            name            = "getMicroTime";
            bOneway         = false;
            cParamInfo[]    = siKernel_getMicroTime_p_system_micro_timeParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo siKernel_getMicroTime_p_system_micro_timeParamInfo {
            name            = "p_system_micro_time";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = SYSUTM_Ptr_TypeInfo.eTypeInfo;
        };

        /*** sSemaphore signature information ****/
        cell nTECSInfo::tSignatureInfo sSemaphoreSignatureInfo {
            name            = "sSemaphore";
            cFunctionInfo[] = sSemaphore_signalFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sSemaphore_waitFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sSemaphore_waitPollingFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sSemaphore_waitTimeoutFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sSemaphore_initializeFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sSemaphore_referFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo sSemaphore_signalFunctionInfo {
            name            = "signal";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sSemaphore_waitFunctionInfo {
            name            = "wait";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sSemaphore_waitPollingFunctionInfo {
            name            = "waitPolling";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sSemaphore_waitTimeoutFunctionInfo {
            name            = "waitTimeout";
            bOneway         = false;
            cParamInfo[]    = sSemaphore_waitTimeout_timeoutParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sSemaphore_waitTimeout_timeoutParamInfo {
            name            = "timeout";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = TMOTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sSemaphore_initializeFunctionInfo {
            name            = "initialize";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sSemaphore_referFunctionInfo {
            name            = "refer";
            bOneway         = false;
            cParamInfo[]    = sSemaphore_refer_pk_semaphore_statusParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sSemaphore_refer_pk_semaphore_statusParamInfo {
            name            = "pk_semaphore_status";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = T_RSEM_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo struct__t_rsem_wtskidVarDeclInfo {
            name            = "wtskid";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_STMEMBER;
            offset          = C_EXP( "OFFSET_OF_struct__t_rsem_wtskid" );
            place           = C_EXP( "PLACE_OF_struct__t_rsem_wtskid" );
            cTypeInfo       = IDTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo struct__t_rsem_semcntVarDeclInfo {
            name            = "semcnt";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_STMEMBER;
            offset          = C_EXP( "OFFSET_OF_struct__t_rsem_semcnt" );
            place           = C_EXP( "PLACE_OF_struct__t_rsem_semcnt" );
            cTypeInfo       = uint_tTypeInfo.eTypeInfo;
        };

        /*** siSemaphore signature information ****/
        cell nTECSInfo::tSignatureInfo siSemaphoreSignatureInfo {
            name            = "siSemaphore";
            cFunctionInfo[] = siSemaphore_signalFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo siSemaphore_signalFunctionInfo {
            name            = "signal";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };

        /*** sEventflag signature information ****/
        cell nTECSInfo::tSignatureInfo sEventflagSignatureInfo {
            name            = "sEventflag";
            cFunctionInfo[] = sEventflag_setFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sEventflag_clearFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sEventflag_waitFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sEventflag_waitPollingFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sEventflag_waitTimeoutFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sEventflag_initializeFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sEventflag_referFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo sEventflag_setFunctionInfo {
            name            = "set";
            bOneway         = false;
            cParamInfo[]    = sEventflag_set_set_patternParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sEventflag_set_set_patternParamInfo {
            name            = "set_pattern";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = FLGPTNTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sEventflag_clearFunctionInfo {
            name            = "clear";
            bOneway         = false;
            cParamInfo[]    = sEventflag_clear_clear_patternParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sEventflag_clear_clear_patternParamInfo {
            name            = "clear_pattern";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = FLGPTNTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sEventflag_waitFunctionInfo {
            name            = "wait";
            bOneway         = false;
            cParamInfo[]    = sEventflag_wait_wait_patternParamInfo.eParamInfo;
            cParamInfo[]    = sEventflag_wait_wait_flag_modeParamInfo.eParamInfo;
            cParamInfo[]    = sEventflag_wait_p_flag_patternParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sEventflag_wait_wait_patternParamInfo {
            name            = "wait_pattern";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = FLGPTNTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sEventflag_wait_wait_flag_modeParamInfo {
            name            = "wait_flag_mode";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = MODETypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sEventflag_wait_p_flag_patternParamInfo {
            name            = "p_flag_pattern";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = FLGPTN_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sEventflag_waitPollingFunctionInfo {
            name            = "waitPolling";
            bOneway         = false;
            cParamInfo[]    = sEventflag_waitPolling_wait_patternParamInfo.eParamInfo;
            cParamInfo[]    = sEventflag_waitPolling_wait_flag_modeParamInfo.eParamInfo;
            cParamInfo[]    = sEventflag_waitPolling_p_flag_patternParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sEventflag_waitPolling_wait_patternParamInfo {
            name            = "wait_pattern";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = FLGPTNTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sEventflag_waitPolling_wait_flag_modeParamInfo {
            name            = "wait_flag_mode";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = MODETypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sEventflag_waitPolling_p_flag_patternParamInfo {
            name            = "p_flag_pattern";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = FLGPTN_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sEventflag_waitTimeoutFunctionInfo {
            name            = "waitTimeout";
            bOneway         = false;
            cParamInfo[]    = sEventflag_waitTimeout_wait_patternParamInfo.eParamInfo;
            cParamInfo[]    = sEventflag_waitTimeout_wait_flag_modeParamInfo.eParamInfo;
            cParamInfo[]    = sEventflag_waitTimeout_p_flag_patternParamInfo.eParamInfo;
            cParamInfo[]    = sEventflag_waitTimeout_timeoutParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sEventflag_waitTimeout_wait_patternParamInfo {
            name            = "wait_pattern";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = FLGPTNTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sEventflag_waitTimeout_wait_flag_modeParamInfo {
            name            = "wait_flag_mode";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = MODETypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sEventflag_waitTimeout_p_flag_patternParamInfo {
            name            = "p_flag_pattern";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = FLGPTN_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sEventflag_waitTimeout_timeoutParamInfo {
            name            = "timeout";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = TMOTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sEventflag_initializeFunctionInfo {
            name            = "initialize";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sEventflag_referFunctionInfo {
            name            = "refer";
            bOneway         = false;
            cParamInfo[]    = sEventflag_refer_pk_eventflag_statusParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sEventflag_refer_pk_eventflag_statusParamInfo {
            name            = "pk_eventflag_status";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = T_RFLG_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo struct__t_rflg_wtskidVarDeclInfo {
            name            = "wtskid";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_STMEMBER;
            offset          = C_EXP( "OFFSET_OF_struct__t_rflg_wtskid" );
            place           = C_EXP( "PLACE_OF_struct__t_rflg_wtskid" );
            cTypeInfo       = IDTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo struct__t_rflg_flgptnVarDeclInfo {
            name            = "flgptn";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_STMEMBER;
            offset          = C_EXP( "OFFSET_OF_struct__t_rflg_flgptn" );
            place           = C_EXP( "PLACE_OF_struct__t_rflg_flgptn" );
            cTypeInfo       = FLGPTNTypeInfo.eTypeInfo;
        };

        /*** siEventflag signature information ****/
        cell nTECSInfo::tSignatureInfo siEventflagSignatureInfo {
            name            = "siEventflag";
            cFunctionInfo[] = siEventflag_setFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo siEventflag_setFunctionInfo {
            name            = "set";
            bOneway         = false;
            cParamInfo[]    = siEventflag_set_set_patternParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo siEventflag_set_set_patternParamInfo {
            name            = "set_pattern";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = FLGPTNTypeInfo.eTypeInfo;
        };

        /*** sDataqueue signature information ****/
        cell nTECSInfo::tSignatureInfo sDataqueueSignatureInfo {
            name            = "sDataqueue";
            cFunctionInfo[] = sDataqueue_sendFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sDataqueue_sendPollingFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sDataqueue_sendTimeoutFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sDataqueue_sendForceFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sDataqueue_receiveFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sDataqueue_receivePollingFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sDataqueue_receiveTimeoutFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sDataqueue_initializeFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = sDataqueue_referFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo sDataqueue_sendFunctionInfo {
            name            = "send";
            bOneway         = false;
            cParamInfo[]    = sDataqueue_send_dataParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sDataqueue_send_dataParamInfo {
            name            = "data";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = intptr_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sDataqueue_sendPollingFunctionInfo {
            name            = "sendPolling";
            bOneway         = false;
            cParamInfo[]    = sDataqueue_sendPolling_dataParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sDataqueue_sendPolling_dataParamInfo {
            name            = "data";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = intptr_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sDataqueue_sendTimeoutFunctionInfo {
            name            = "sendTimeout";
            bOneway         = false;
            cParamInfo[]    = sDataqueue_sendTimeout_dataParamInfo.eParamInfo;
            cParamInfo[]    = sDataqueue_sendTimeout_timeoutParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sDataqueue_sendTimeout_dataParamInfo {
            name            = "data";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = intptr_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sDataqueue_sendTimeout_timeoutParamInfo {
            name            = "timeout";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = TMOTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sDataqueue_sendForceFunctionInfo {
            name            = "sendForce";
            bOneway         = false;
            cParamInfo[]    = sDataqueue_sendForce_dataParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sDataqueue_sendForce_dataParamInfo {
            name            = "data";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = intptr_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sDataqueue_receiveFunctionInfo {
            name            = "receive";
            bOneway         = false;
            cParamInfo[]    = sDataqueue_receive_p_dataParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sDataqueue_receive_p_dataParamInfo {
            name            = "p_data";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = intptr_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sDataqueue_receivePollingFunctionInfo {
            name            = "receivePolling";
            bOneway         = false;
            cParamInfo[]    = sDataqueue_receivePolling_p_dataParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sDataqueue_receivePolling_p_dataParamInfo {
            name            = "p_data";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = intptr_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sDataqueue_receiveTimeoutFunctionInfo {
            name            = "receiveTimeout";
            bOneway         = false;
            cParamInfo[]    = sDataqueue_receiveTimeout_p_dataParamInfo.eParamInfo;
            cParamInfo[]    = sDataqueue_receiveTimeout_timeoutParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sDataqueue_receiveTimeout_p_dataParamInfo {
            name            = "p_data";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = intptr_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sDataqueue_receiveTimeout_timeoutParamInfo {
            name            = "timeout";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = TMOTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sDataqueue_initializeFunctionInfo {
            name            = "initialize";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo sDataqueue_referFunctionInfo {
            name            = "refer";
            bOneway         = false;
            cParamInfo[]    = sDataqueue_refer_pk_dataqueue_statusParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sDataqueue_refer_pk_dataqueue_statusParamInfo {
            name            = "pk_dataqueue_status";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = T_RDTQ_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo struct__t_rdtq_stskidVarDeclInfo {
            name            = "stskid";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_STMEMBER;
            offset          = C_EXP( "OFFSET_OF_struct__t_rdtq_stskid" );
            place           = C_EXP( "PLACE_OF_struct__t_rdtq_stskid" );
            cTypeInfo       = IDTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo struct__t_rdtq_rtskidVarDeclInfo {
            name            = "rtskid";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_STMEMBER;
            offset          = C_EXP( "OFFSET_OF_struct__t_rdtq_rtskid" );
            place           = C_EXP( "PLACE_OF_struct__t_rdtq_rtskid" );
            cTypeInfo       = IDTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo struct__t_rdtq_sdtqcntVarDeclInfo {
            name            = "sdtqcnt";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_STMEMBER;
            offset          = C_EXP( "OFFSET_OF_struct__t_rdtq_sdtqcnt" );
            place           = C_EXP( "PLACE_OF_struct__t_rdtq_sdtqcnt" );
            cTypeInfo       = uint_tTypeInfo.eTypeInfo;
        };

        /*** siDataqueue signature information ****/
        cell nTECSInfo::tSignatureInfo siDataqueueSignatureInfo {
            name            = "siDataqueue";
            cFunctionInfo[] = siDataqueue_sendPollingFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = siDataqueue_sendForceFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo siDataqueue_sendPollingFunctionInfo {
            name            = "sendPolling";
            bOneway         = false;
            cParamInfo[]    = siDataqueue_sendPolling_dataParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo siDataqueue_sendPolling_dataParamInfo {
            name            = "data";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = intptr_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo siDataqueue_sendForceFunctionInfo {
            name            = "sendForce";
            bOneway         = false;
            cParamInfo[]    = siDataqueue_sendForce_dataParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo siDataqueue_sendForce_dataParamInfo {
            name            = "data";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = intptr_tTypeInfo.eTypeInfo;
        };

        /*** sPutString signature information ****/
        cell nTECSInfo::tSignatureInfo sPutStringSignatureInfo {
            name            = "sPutString";
            cFunctionInfo[] = sPutString_putStringFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo sPutString_putStringFunctionInfo {
            name            = "putString";
            bOneway         = false;
            cParamInfo[]    = sPutString_putString_stringParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo sPutString_putString_stringParamInfo {
            name            = "string";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tCelltypeInfo tTaskCelltypeInfo {
            name             = "tTask";
            b_singleton      = false;
            b_IDX_is_ID_act  = C_EXP( "tTask__IDX_is_ID_act" );
            sizeOfCB         = C_EXP( "tTask__sizeOfCB" );
            sizeOfINIB       = C_EXP( "tTask__sizeOfINIB" );
            n_cellInLinkUnit = C_EXP( "tTask__NCELLINLINKUNIT" );
            n_cellInSystem   = 1;
            cEntryInfo[]    = tTask_eTaskEntryInfo.eEntryInfo;
            cCallInfo[]     = tTask_cTaskBodyCallInfo.eCallInfo;
            cCallInfo[]     = tTask_cExceptionBodyCallInfo.eCallInfo;
            cAttrInfo[]     = tTask_attributeVarDeclInfo.eVarDeclInfo;
            cAttrInfo[]     = tTask_priorityVarDeclInfo.eVarDeclInfo;
            cAttrInfo[]     = tTask_stackSizeVarDeclInfo.eVarDeclInfo;
            cAttrInfo[]     = tTask_nameVarDeclInfo.eVarDeclInfo;
            cVarInfo[]      = tTask_my_threadVarDeclInfo.eVarDeclInfo;
            cVarInfo[]      = tTask_my_condVarDeclInfo.eVarDeclInfo;
            cVarInfo[]      = tTask_my_mutexVarDeclInfo.eVarDeclInfo;
            cVarInfo[]      = tTask_stateVarDeclInfo.eVarDeclInfo;
        };
        cell nTECSInfo::tEntryInfo tTask_eTaskEntryInfo{
            name            = "eTask";
            cSignatureInfo  = sTaskSignatureInfo.eSignatureInfo;
            b_inline        = true;
            array_size      = C_EXP( "tTask_eTask__array_size" );
        };
        cell nTECSInfo::tCallInfo tTask_cTaskBodyCallInfo{
            name            = "cTaskBody";
            cSignatureInfo  = sTaskBodySignatureInfo.eSignatureInfo;
            offset            = C_EXP( "tTask_cTaskBody__offset" );
            array_size        = C_EXP( "tTask_cTaskBody__array_size" );
            b_optional        = false;
            b_omit            = false;
            b_dynamic         = false;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "tTask_cTaskBody__place" );
            b_VMT_useless     = C_EXP( "tTask_cTaskBody__b_VMT_useless" );
            b_skelton_useless = C_EXP( "tTask_cTaskBody__b_skelton_useless" );
            b_cell_unique     = C_EXP( "tTask_cTaskBody__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo tTask_cExceptionBodyCallInfo{
            name            = "cExceptionBody";
            cSignatureInfo  = sTaskExceptionBodySignatureInfo.eSignatureInfo;
            offset            = C_EXP( "tTask_cExceptionBody__offset" );
            array_size        = C_EXP( "tTask_cExceptionBody__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = false;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "tTask_cExceptionBody__place" );
            b_VMT_useless     = C_EXP( "tTask_cExceptionBody__b_VMT_useless" );
            b_skelton_useless = C_EXP( "tTask_cExceptionBody__b_skelton_useless" );
            b_cell_unique     = C_EXP( "tTask_cExceptionBody__b_cell_unique" );

        };
        cell nTECSInfo::tVarDeclInfo tTask_attributeVarDeclInfo {
            name            = "attribute";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_ATTR;
            offset          = C_EXP( "OFFSET_OF_tTask_attribute" );
            place           = C_EXP( "PLACE_OF_tTask_attribute" );
            cTypeInfo       = ATRTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo tTask_priorityVarDeclInfo {
            name            = "priority";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_ATTR;
            offset          = C_EXP( "OFFSET_OF_tTask_priority" );
            place           = C_EXP( "PLACE_OF_tTask_priority" );
            cTypeInfo       = PRITypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo tTask_stackSizeVarDeclInfo {
            name            = "stackSize";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_ATTR;
            offset          = C_EXP( "OFFSET_OF_tTask_stackSize" );
            place           = C_EXP( "PLACE_OF_tTask_stackSize" );
            cTypeInfo       = size_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo tTask_nameVarDeclInfo {
            name            = "name";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_ATTR;
            offset          = C_EXP( "OFFSET_OF_tTask_name" );
            place           = C_EXP( "PLACE_OF_tTask_name" );
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo tTask_my_threadVarDeclInfo {
            name            = "my_thread";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_VAR;
            offset          = C_EXP( "OFFSET_OF_tTask_my_thread" );
            place           = C_EXP( "PLACE_OF_tTask_my_thread" );
            cTypeInfo       = pthread_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo tTask_my_condVarDeclInfo {
            name            = "my_cond";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_VAR;
            offset          = C_EXP( "OFFSET_OF_tTask_my_cond" );
            place           = C_EXP( "PLACE_OF_tTask_my_cond" );
            cTypeInfo       = pthread_cond_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo tTask_my_mutexVarDeclInfo {
            name            = "my_mutex";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_VAR;
            offset          = C_EXP( "OFFSET_OF_tTask_my_mutex" );
            place           = C_EXP( "PLACE_OF_tTask_my_mutex" );
            cTypeInfo       = pthread_mutex_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo tTask_stateVarDeclInfo {
            name            = "state";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_VAR;
            offset          = C_EXP( "OFFSET_OF_tTask_state" );
            place           = C_EXP( "PLACE_OF_tTask_state" );
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tCelltypeInfo tPutStringStdioCelltypeInfo {
            name             = "tPutStringStdio";
            b_singleton      = false;
            b_IDX_is_ID_act  = C_EXP( "tPutStringStdio__IDX_is_ID_act" );
            sizeOfCB         = C_EXP( "tPutStringStdio__sizeOfCB" );
            sizeOfINIB       = C_EXP( "tPutStringStdio__sizeOfINIB" );
            n_cellInLinkUnit = C_EXP( "tPutStringStdio__NCELLINLINKUNIT" );
            n_cellInSystem   = 1;
            cEntryInfo[]    = tPutStringStdio_ePutStringEntryInfo.eEntryInfo;
        };
        cell nTECSInfo::tEntryInfo tPutStringStdio_ePutStringEntryInfo{
            name            = "ePutString";
            cSignatureInfo  = sPutStringSignatureInfo.eSignatureInfo;
            b_inline        = false;
            array_size      = C_EXP( "tPutStringStdio_ePutString__array_size" );
        };
        cell nTECSInfo::tCelltypeInfo tHelloWorldCelltypeInfo {
            name             = "tHelloWorld";
            b_singleton      = false;
            b_IDX_is_ID_act  = C_EXP( "tHelloWorld__IDX_is_ID_act" );
            sizeOfCB         = C_EXP( "tHelloWorld__sizeOfCB" );
            sizeOfINIB       = C_EXP( "tHelloWorld__sizeOfINIB" );
            n_cellInLinkUnit = C_EXP( "tHelloWorld__NCELLINLINKUNIT" );
            n_cellInSystem   = 1;
            cEntryInfo[]    = tHelloWorld_eMainEntryInfo.eEntryInfo;
            cCallInfo[]     = tHelloWorld_cPutStringCallInfo.eCallInfo;
            cAttrInfo[]     = tHelloWorld_messageVarDeclInfo.eVarDeclInfo;
        };
        cell nTECSInfo::tEntryInfo tHelloWorld_eMainEntryInfo{
            name            = "eMain";
            cSignatureInfo  = sTaskBodySignatureInfo.eSignatureInfo;
            b_inline        = false;
            array_size      = C_EXP( "tHelloWorld_eMain__array_size" );
        };
        cell nTECSInfo::tCallInfo tHelloWorld_cPutStringCallInfo{
            name            = "cPutString";
            cSignatureInfo  = sPutStringSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "tHelloWorld_cPutString__offset" );
            array_size        = C_EXP( "tHelloWorld_cPutString__array_size" );
            b_optional        = false;
            b_omit            = false;
            b_dynamic         = false;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "tHelloWorld_cPutString__place" );
            b_VMT_useless     = C_EXP( "tHelloWorld_cPutString__b_VMT_useless" );
            b_skelton_useless = C_EXP( "tHelloWorld_cPutString__b_skelton_useless" );
            b_cell_unique     = C_EXP( "tHelloWorld_cPutString__b_cell_unique" );

        };
        cell nTECSInfo::tVarDeclInfo tHelloWorld_messageVarDeclInfo {
            name            = "message";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_ATTR;
            offset          = C_EXP( "OFFSET_OF_tHelloWorld_message" );
            place           = C_EXP( "PLACE_OF_tHelloWorld_message" );
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tCelltypeInfo tTaskMainCelltypeInfo {
            name             = "tTaskMain";
            b_singleton      = false;
            b_IDX_is_ID_act  = C_EXP( "tTaskMain__IDX_is_ID_act" );
            sizeOfCB         = C_EXP( "tTaskMain__sizeOfCB" );
            sizeOfINIB       = C_EXP( "tTaskMain__sizeOfINIB" );
            n_cellInLinkUnit = C_EXP( "tTaskMain__NCELLINLINKUNIT" );
            n_cellInSystem   = 1;
            cEntryInfo[]    = tTaskMain_eBodyEntryInfo.eEntryInfo;
            cCallInfo[]     = tTaskMain_cAccessorCallInfo.eCallInfo;
            cAttrInfo[]     = tTaskMain_NAME_LENVarDeclInfo.eVarDeclInfo;
            cVarInfo[]      = tTaskMain_nameVarDeclInfo.eVarDeclInfo;
            cVarInfo[]      = tTaskMain_name2VarDeclInfo.eVarDeclInfo;
        };
        cell nTECSInfo::tEntryInfo tTaskMain_eBodyEntryInfo{
            name            = "eBody";
            cSignatureInfo  = sTaskBodySignatureInfo.eSignatureInfo;
            b_inline        = false;
            array_size      = C_EXP( "tTaskMain_eBody__array_size" );
        };
        cell nTECSInfo::tCallInfo tTaskMain_cAccessorCallInfo{
            name            = "cAccessor";
            cSignatureInfo  = nTECSInfo_sAccessorSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "tTaskMain_cAccessor__offset" );
            array_size        = C_EXP( "tTaskMain_cAccessor__array_size" );
            b_optional        = false;
            b_omit            = false;
            b_dynamic         = false;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "tTaskMain_cAccessor__place" );
            b_VMT_useless     = C_EXP( "tTaskMain_cAccessor__b_VMT_useless" );
            b_skelton_useless = C_EXP( "tTaskMain_cAccessor__b_skelton_useless" );
            b_cell_unique     = C_EXP( "tTaskMain_cAccessor__b_cell_unique" );

        };
        cell nTECSInfo::tVarDeclInfo tTaskMain_NAME_LENVarDeclInfo {
            name            = "NAME_LEN";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_ATTR;
            offset          = C_EXP( "OFFSET_OF_tTaskMain_NAME_LEN" );
            place           = C_EXP( "PLACE_OF_tTaskMain_NAME_LEN" );
            cTypeInfo       = int16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo tTaskMain_nameVarDeclInfo {
            name            = "name";
            sizeIsExpr      = "mikan";
            declType        = DECLTYPE_VAR;
            offset          = C_EXP( "OFFSET_OF_tTaskMain_name" );
            place           = C_EXP( "PLACE_OF_tTaskMain_name" );
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo tTaskMain_name2VarDeclInfo {
            name            = "name2";
            sizeIsExpr      = "mikan";
            declType        = DECLTYPE_VAR;
            offset          = C_EXP( "OFFSET_OF_tTaskMain_name2" );
            place           = C_EXP( "PLACE_OF_tTaskMain_name2" );
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };

        /*** ::nTECSInfo namespace information cell ***/
        cell nTECSInfo::tNamespaceInfo nTECSInfoNamespaceInfo{
            name = "nTECSInfo";

            /* SIGNATURE info */
            cSignatureInfo[] = nTECSInfo_sTypeInfoSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = nTECSInfo_sVarDeclInfoSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = nTECSInfo_sParamInfoSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = nTECSInfo_sFunctionInfoSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = nTECSInfo_sSignatureInfoSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = nTECSInfo_sCallInfoSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = nTECSInfo_sEntryInfoSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = nTECSInfo_sCelltypeInfoSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = nTECSInfo_sCellInfoSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = nTECSInfo_sRawEntryDescriptorInfoSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = nTECSInfo_sNamespaceInfoSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = nTECSInfo_sRegionInfoSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = nTECSInfo_sTECSInfoSignatureInfo.eSignatureInfo;
            cSignatureInfo[] = nTECSInfo_sAccessorSignatureInfo.eSignatureInfo;

            /* CELLTYPE info */
            cCelltypeInfo[] = nTECSInfo_tTECSInfoCelltypeInfo.eCelltypeInfo;
            cCelltypeInfo[] = nTECSInfo_tTECSInfoAccessorCelltypeInfo.eCelltypeInfo;
        };   /* cell nTECSInfo::tNamespaceInfo nTECSInfoNamespaceInfo */

        /*** nTECSInfo_sTypeInfo signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sTypeInfoSignatureInfo {
            name            = "sTypeInfo";
            cFunctionInfo[] = nTECSInfo_sTypeInfo_getNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sTypeInfo_getNameLengthFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sTypeInfo_getSizeFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sTypeInfo_getKindFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sTypeInfo_getNTypeFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sTypeInfo_getTypeInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sTypeInfo_getNMemberFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sTypeInfo_getMemberInfoFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTypeInfo_getNameFunctionInfo {
            name            = "getName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sTypeInfo_getName_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sTypeInfo_getName_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTypeInfo_getName_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTypeInfo_getName_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTypeInfo_getNameLengthFunctionInfo {
            name            = "getNameLength";
            bOneway         = false;
            cReturnTypeInfo = uint16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTypeInfo_getSizeFunctionInfo {
            name            = "getSize";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTypeInfo_getKindFunctionInfo {
            name            = "getKind";
            bOneway         = false;
            cReturnTypeInfo = int8_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTypeInfo_getNTypeFunctionInfo {
            name            = "getNType";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTypeInfo_getTypeInfoFunctionInfo {
            name            = "getTypeInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sTypeInfo_getTypeInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTypeInfo_getTypeInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sTypeInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTypeInfo_getNMemberFunctionInfo {
            name            = "getNMember";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTypeInfo_getMemberInfoFunctionInfo {
            name            = "getMemberInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sTypeInfo_getMemberInfo_ithParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sTypeInfo_getMemberInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTypeInfo_getMemberInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTypeInfo_getMemberInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sVarDeclInfo_Ptr_TypeInfo.eTypeInfo;
        };

        /*** nTECSInfo_sVarDeclInfo signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sVarDeclInfoSignatureInfo {
            name            = "sVarDeclInfo";
            cFunctionInfo[] = nTECSInfo_sVarDeclInfo_getNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sVarDeclInfo_getNameLengthFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sVarDeclInfo_getLocationInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sVarDeclInfo_getTypeInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sVarDeclInfo_getSizeIsExprFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sVarDeclInfo_getSizeIsFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sVarDeclInfo_getNameFunctionInfo {
            name            = "getName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sVarDeclInfo_getName_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sVarDeclInfo_getName_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sVarDeclInfo_getName_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sVarDeclInfo_getName_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sVarDeclInfo_getNameLengthFunctionInfo {
            name            = "getNameLength";
            bOneway         = false;
            cReturnTypeInfo = uint16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sVarDeclInfo_getLocationInfoFunctionInfo {
            name            = "getLocationInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sVarDeclInfo_getLocationInfo_offsetParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sVarDeclInfo_getLocationInfo_placeParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sVarDeclInfo_getLocationInfo_offsetParamInfo {
            name            = "offset";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sVarDeclInfo_getLocationInfo_placeParamInfo {
            name            = "place";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int8_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sVarDeclInfo_getTypeInfoFunctionInfo {
            name            = "getTypeInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sVarDeclInfo_getTypeInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sVarDeclInfo_getTypeInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sTypeInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sVarDeclInfo_getSizeIsExprFunctionInfo {
            name            = "getSizeIsExpr";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sVarDeclInfo_getSizeIsExpr_expr_strParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sVarDeclInfo_getSizeIsExpr_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sVarDeclInfo_getSizeIsExpr_expr_strParamInfo {
            name            = "expr_str";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sVarDeclInfo_getSizeIsExpr_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sVarDeclInfo_getSizeIsFunctionInfo {
            name            = "getSizeIs";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sVarDeclInfo_getSizeIs_sizeParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sVarDeclInfo_getSizeIs_p_cbParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sVarDeclInfo_getSizeIs_sizeParamInfo {
            name            = "size";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sVarDeclInfo_getSizeIs_p_cbParamInfo {
            name            = "p_cb";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = const__void_Ptr_TypeInfo.eTypeInfo;
        };

        /*** nTECSInfo_sParamInfo signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sParamInfoSignatureInfo {
            name            = "sParamInfo";
            cFunctionInfo[] = nTECSInfo_sParamInfo_getNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sParamInfo_getNameLengthFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sParamInfo_getTypeInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sParamInfo_getDirFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sParamInfo_getNameFunctionInfo {
            name            = "getName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sParamInfo_getName_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sParamInfo_getName_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sParamInfo_getName_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sParamInfo_getName_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sParamInfo_getNameLengthFunctionInfo {
            name            = "getNameLength";
            bOneway         = false;
            cReturnTypeInfo = uint16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sParamInfo_getTypeInfoFunctionInfo {
            name            = "getTypeInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sParamInfo_getTypeInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sParamInfo_getTypeInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sTypeInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sParamInfo_getDirFunctionInfo {
            name            = "getDir";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sParamInfo_getDir_dirParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sParamInfo_getDir_dirParamInfo {
            name            = "dir";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int8_t_Ptr_TypeInfo.eTypeInfo;
        };

        /*** nTECSInfo_sFunctionInfo signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sFunctionInfoSignatureInfo {
            name            = "sFunctionInfo";
            cFunctionInfo[] = nTECSInfo_sFunctionInfo_getNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sFunctionInfo_getNameLengthFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sFunctionInfo_getReturnTypeInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sFunctionInfo_getNParamFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sFunctionInfo_getParamInfoFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sFunctionInfo_getNameFunctionInfo {
            name            = "getName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sFunctionInfo_getName_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sFunctionInfo_getName_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sFunctionInfo_getName_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sFunctionInfo_getName_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sFunctionInfo_getNameLengthFunctionInfo {
            name            = "getNameLength";
            bOneway         = false;
            cReturnTypeInfo = uint16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sFunctionInfo_getReturnTypeInfoFunctionInfo {
            name            = "getReturnTypeInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sFunctionInfo_getReturnTypeInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sFunctionInfo_getReturnTypeInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sTypeInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sFunctionInfo_getNParamFunctionInfo {
            name            = "getNParam";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sFunctionInfo_getParamInfoFunctionInfo {
            name            = "getParamInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sFunctionInfo_getParamInfo_ithParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sFunctionInfo_getParamInfo_paramParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sFunctionInfo_getParamInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sFunctionInfo_getParamInfo_paramParamInfo {
            name            = "param";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sParamInfo_Ptr_TypeInfo.eTypeInfo;
        };

        /*** nTECSInfo_sSignatureInfo signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sSignatureInfoSignatureInfo {
            name            = "sSignatureInfo";
            cFunctionInfo[] = nTECSInfo_sSignatureInfo_getNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sSignatureInfo_getNameLengthFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sSignatureInfo_getNFunctionFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sSignatureInfo_getFunctionInfoFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sSignatureInfo_getNameFunctionInfo {
            name            = "getName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sSignatureInfo_getName_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sSignatureInfo_getName_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sSignatureInfo_getName_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sSignatureInfo_getName_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sSignatureInfo_getNameLengthFunctionInfo {
            name            = "getNameLength";
            bOneway         = false;
            cReturnTypeInfo = uint16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sSignatureInfo_getNFunctionFunctionInfo {
            name            = "getNFunction";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sSignatureInfo_getFunctionInfoFunctionInfo {
            name            = "getFunctionInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sSignatureInfo_getFunctionInfo_ithParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sSignatureInfo_getFunctionInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sSignatureInfo_getFunctionInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sSignatureInfo_getFunctionInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sFunctionInfo_Ptr_TypeInfo.eTypeInfo;
        };

        /*** nTECSInfo_sCallInfo signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sCallInfoSignatureInfo {
            name            = "sCallInfo";
            cFunctionInfo[] = nTECSInfo_sCallInfo_getNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCallInfo_getNameLengthFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCallInfo_getSignatureInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCallInfo_getArraySizeFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCallInfo_getSpecifierInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCallInfo_getInternalInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCallInfo_getLocationInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCallInfo_getOptimizeInfoFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCallInfo_getNameFunctionInfo {
            name            = "getName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCallInfo_getName_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCallInfo_getName_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getName_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getName_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCallInfo_getNameLengthFunctionInfo {
            name            = "getNameLength";
            bOneway         = false;
            cReturnTypeInfo = uint16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCallInfo_getSignatureInfoFunctionInfo {
            name            = "getSignatureInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCallInfo_getSignatureInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getSignatureInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sSignatureInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCallInfo_getArraySizeFunctionInfo {
            name            = "getArraySize";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCallInfo_getSpecifierInfoFunctionInfo {
            name            = "getSpecifierInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCallInfo_getSpecifierInfo_b_optionalParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCallInfo_getSpecifierInfo_b_dynamicParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCallInfo_getSpecifierInfo_b_ref_descParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCallInfo_getSpecifierInfo_b_omitParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getSpecifierInfo_b_optionalParamInfo {
            name            = "b_optional";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getSpecifierInfo_b_dynamicParamInfo {
            name            = "b_dynamic";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getSpecifierInfo_b_ref_descParamInfo {
            name            = "b_ref_desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getSpecifierInfo_b_omitParamInfo {
            name            = "b_omit";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCallInfo_getInternalInfoFunctionInfo {
            name            = "getInternalInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCallInfo_getInternalInfo_b_allocator_portParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCallInfo_getInternalInfo_b_require_portParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getInternalInfo_b_allocator_portParamInfo {
            name            = "b_allocator_port";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getInternalInfo_b_require_portParamInfo {
            name            = "b_require_port";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCallInfo_getLocationInfoFunctionInfo {
            name            = "getLocationInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCallInfo_getLocationInfo_offsetParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCallInfo_getLocationInfo_placeParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getLocationInfo_offsetParamInfo {
            name            = "offset";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getLocationInfo_placeParamInfo {
            name            = "place";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int8_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCallInfo_getOptimizeInfoFunctionInfo {
            name            = "getOptimizeInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCallInfo_getOptimizeInfo_b_VMT_uselessParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCallInfo_getOptimizeInfo_b_skelton_uselessParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCallInfo_getOptimizeInfo_b_cell_uniqueParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getOptimizeInfo_b_VMT_uselessParamInfo {
            name            = "b_VMT_useless";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getOptimizeInfo_b_skelton_uselessParamInfo {
            name            = "b_skelton_useless";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCallInfo_getOptimizeInfo_b_cell_uniqueParamInfo {
            name            = "b_cell_unique";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };

        /*** nTECSInfo_sEntryInfo signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sEntryInfoSignatureInfo {
            name            = "sEntryInfo";
            cFunctionInfo[] = nTECSInfo_sEntryInfo_getNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sEntryInfo_getNameLengthFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sEntryInfo_getSignatureInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sEntryInfo_getArraySizeFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sEntryInfo_isInlineFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sEntryInfo_getNameFunctionInfo {
            name            = "getName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sEntryInfo_getName_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sEntryInfo_getName_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sEntryInfo_getName_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sEntryInfo_getName_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sEntryInfo_getNameLengthFunctionInfo {
            name            = "getNameLength";
            bOneway         = false;
            cReturnTypeInfo = uint16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sEntryInfo_getSignatureInfoFunctionInfo {
            name            = "getSignatureInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sEntryInfo_getSignatureInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sEntryInfo_getSignatureInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sSignatureInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sEntryInfo_getArraySizeFunctionInfo {
            name            = "getArraySize";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sEntryInfo_isInlineFunctionInfo {
            name            = "isInline";
            bOneway         = false;
            cReturnTypeInfo = bool_tTypeInfo.eTypeInfo;
        };

        /*** nTECSInfo_sCelltypeInfo signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sCelltypeInfoSignatureInfo {
            name            = "sCelltypeInfo";
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_getNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_getNameLengthFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_getNAttrFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_getAttrInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_getNVarFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_getVarInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_getNCallFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_getCallInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_getNEntryFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_getEntryInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_isSingletonFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_isIDX_is_IDFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_sizeOfCBFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCelltypeInfo_sizeOfINIBFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_getNameFunctionInfo {
            name            = "getName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCelltypeInfo_getName_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCelltypeInfo_getName_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCelltypeInfo_getName_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCelltypeInfo_getName_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_getNameLengthFunctionInfo {
            name            = "getNameLength";
            bOneway         = false;
            cReturnTypeInfo = uint16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_getNAttrFunctionInfo {
            name            = "getNAttr";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_getAttrInfoFunctionInfo {
            name            = "getAttrInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCelltypeInfo_getAttrInfo_ithParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCelltypeInfo_getAttrInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCelltypeInfo_getAttrInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCelltypeInfo_getAttrInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sVarDeclInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_getNVarFunctionInfo {
            name            = "getNVar";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_getVarInfoFunctionInfo {
            name            = "getVarInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCelltypeInfo_getVarInfo_ithParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCelltypeInfo_getVarInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCelltypeInfo_getVarInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCelltypeInfo_getVarInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sVarDeclInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_getNCallFunctionInfo {
            name            = "getNCall";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_getCallInfoFunctionInfo {
            name            = "getCallInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCelltypeInfo_getCallInfo_ithParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCelltypeInfo_getCallInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCelltypeInfo_getCallInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCelltypeInfo_getCallInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sCallInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_getNEntryFunctionInfo {
            name            = "getNEntry";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_getEntryInfoFunctionInfo {
            name            = "getEntryInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCelltypeInfo_getEntryInfo_ithParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCelltypeInfo_getEntryInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCelltypeInfo_getEntryInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCelltypeInfo_getEntryInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sEntryInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_isSingletonFunctionInfo {
            name            = "isSingleton";
            bOneway         = false;
            cReturnTypeInfo = bool_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_isIDX_is_IDFunctionInfo {
            name            = "isIDX_is_ID";
            bOneway         = false;
            cReturnTypeInfo = bool_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_sizeOfCBFunctionInfo {
            name            = "sizeOfCB";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCelltypeInfo_sizeOfINIBFunctionInfo {
            name            = "sizeOfINIB";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };

        /*** nTECSInfo_sCellInfo signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sCellInfoSignatureInfo {
            name            = "sCellInfo";
            cFunctionInfo[] = nTECSInfo_sCellInfo_getNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCellInfo_getNameLengthFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCellInfo_getNRawEntryDescriptorInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCellInfo_getRawEntryDescriptorInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCellInfo_getCelltypeInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCellInfo_getCBPFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sCellInfo_getINIBPFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCellInfo_getNameFunctionInfo {
            name            = "getName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCellInfo_getName_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCellInfo_getName_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCellInfo_getName_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCellInfo_getName_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCellInfo_getNameLengthFunctionInfo {
            name            = "getNameLength";
            bOneway         = false;
            cReturnTypeInfo = uint16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCellInfo_getNRawEntryDescriptorInfoFunctionInfo {
            name            = "getNRawEntryDescriptorInfo";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCellInfo_getRawEntryDescriptorInfoFunctionInfo {
            name            = "getRawEntryDescriptorInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCellInfo_getRawEntryDescriptorInfo_indexParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sCellInfo_getRawEntryDescriptorInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCellInfo_getRawEntryDescriptorInfo_indexParamInfo {
            name            = "index";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCellInfo_getRawEntryDescriptorInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sRawEntryDescriptorInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCellInfo_getCelltypeInfoFunctionInfo {
            name            = "getCelltypeInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCellInfo_getCelltypeInfo_descParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCellInfo_getCelltypeInfo_descParamInfo {
            name            = "desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sCelltypeInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCellInfo_getCBPFunctionInfo {
            name            = "getCBP";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCellInfo_getCBP_cbpParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCellInfo_getCBP_cbpParamInfo {
            name            = "cbp";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = void_Ptr__Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sCellInfo_getINIBPFunctionInfo {
            name            = "getINIBP";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sCellInfo_getINIBP_inibpParamInfo.eParamInfo;
            cReturnTypeInfo = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sCellInfo_getINIBP_inibpParamInfo {
            name            = "inibp";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = void_Ptr__Ptr_TypeInfo.eTypeInfo;
        };

        /*** nTECSInfo_sRawEntryDescriptorInfo signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sRawEntryDescriptorInfoSignatureInfo {
            name            = "sRawEntryDescriptorInfo";
            cFunctionInfo[] = nTECSInfo_sRawEntryDescriptorInfo_getNRawEntryDescriptorInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sRawEntryDescriptorInfo_getRawDescriptorFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sRawEntryDescriptorInfo_getNRawEntryDescriptorInfoFunctionInfo {
            name            = "getNRawEntryDescriptorInfo";
            bOneway         = false;
            cReturnTypeInfo = uint16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sRawEntryDescriptorInfo_getRawDescriptorFunctionInfo {
            name            = "getRawDescriptor";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sRawEntryDescriptorInfo_getRawDescriptor_subscParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sRawEntryDescriptorInfo_getRawDescriptor_rawDescParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sRawEntryDescriptorInfo_getRawDescriptor_subscParamInfo {
            name            = "subsc";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sRawEntryDescriptorInfo_getRawDescriptor_rawDescParamInfo {
            name            = "rawDesc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = void_Ptr__Ptr_TypeInfo.eTypeInfo;
        };

        /*** nTECSInfo_sNamespaceInfo signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sNamespaceInfoSignatureInfo {
            name            = "sNamespaceInfo";
            cFunctionInfo[] = nTECSInfo_sNamespaceInfo_getNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sNamespaceInfo_getNameLengthFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sNamespaceInfo_getNNamespaceFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sNamespaceInfo_getNamespaceInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sNamespaceInfo_getNSignatureFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sNamespaceInfo_getSignatureInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sNamespaceInfo_getNCelltypeFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sNamespaceInfo_getCelltypeInfoFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sNamespaceInfo_getNameFunctionInfo {
            name            = "getName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sNamespaceInfo_getName_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sNamespaceInfo_getName_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sNamespaceInfo_getName_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sNamespaceInfo_getName_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sNamespaceInfo_getNameLengthFunctionInfo {
            name            = "getNameLength";
            bOneway         = false;
            cReturnTypeInfo = uint16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sNamespaceInfo_getNNamespaceFunctionInfo {
            name            = "getNNamespace";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sNamespaceInfo_getNamespaceInfoFunctionInfo {
            name            = "getNamespaceInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sNamespaceInfo_getNamespaceInfo_ithParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sNamespaceInfo_getNamespaceInfo_desParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sNamespaceInfo_getNamespaceInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sNamespaceInfo_getNamespaceInfo_desParamInfo {
            name            = "des";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sNamespaceInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sNamespaceInfo_getNSignatureFunctionInfo {
            name            = "getNSignature";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sNamespaceInfo_getSignatureInfoFunctionInfo {
            name            = "getSignatureInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sNamespaceInfo_getSignatureInfo_ithParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sNamespaceInfo_getSignatureInfo_desParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sNamespaceInfo_getSignatureInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sNamespaceInfo_getSignatureInfo_desParamInfo {
            name            = "des";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sSignatureInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sNamespaceInfo_getNCelltypeFunctionInfo {
            name            = "getNCelltype";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sNamespaceInfo_getCelltypeInfoFunctionInfo {
            name            = "getCelltypeInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sNamespaceInfo_getCelltypeInfo_ithParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sNamespaceInfo_getCelltypeInfo_desParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sNamespaceInfo_getCelltypeInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sNamespaceInfo_getCelltypeInfo_desParamInfo {
            name            = "des";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sCelltypeInfo_Ptr_TypeInfo.eTypeInfo;
        };

        /*** nTECSInfo_sRegionInfo signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sRegionInfoSignatureInfo {
            name            = "sRegionInfo";
            cFunctionInfo[] = nTECSInfo_sRegionInfo_getNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sRegionInfo_getNameLengthFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sRegionInfo_getNCellFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sRegionInfo_getCellInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sRegionInfo_getNRegionFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sRegionInfo_getRegionInfoFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sRegionInfo_getNameFunctionInfo {
            name            = "getName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sRegionInfo_getName_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sRegionInfo_getName_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sRegionInfo_getName_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sRegionInfo_getName_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sRegionInfo_getNameLengthFunctionInfo {
            name            = "getNameLength";
            bOneway         = false;
            cReturnTypeInfo = uint16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sRegionInfo_getNCellFunctionInfo {
            name            = "getNCell";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sRegionInfo_getCellInfoFunctionInfo {
            name            = "getCellInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sRegionInfo_getCellInfo_ithParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sRegionInfo_getCellInfo_desParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sRegionInfo_getCellInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sRegionInfo_getCellInfo_desParamInfo {
            name            = "des";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sCellInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sRegionInfo_getNRegionFunctionInfo {
            name            = "getNRegion";
            bOneway         = false;
            cReturnTypeInfo = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sRegionInfo_getRegionInfoFunctionInfo {
            name            = "getRegionInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sRegionInfo_getRegionInfo_ithParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sRegionInfo_getRegionInfo_desParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sRegionInfo_getRegionInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sRegionInfo_getRegionInfo_desParamInfo {
            name            = "des";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sRegionInfo_Ptr_TypeInfo.eTypeInfo;
        };

        /*** nTECSInfo_sTECSInfo signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sTECSInfoSignatureInfo {
            name            = "sTECSInfo";
            cFunctionInfo[] = nTECSInfo_sTECSInfo_findNamespaceFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sTECSInfo_findRegionFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sTECSInfo_findSignatureFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sTECSInfo_findCelltypeFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sTECSInfo_findCellFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sTECSInfo_findRawEntryDescriptorFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sTECSInfo_findRawEntryDescriptor_unsafeFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTECSInfo_findNamespaceFunctionInfo {
            name            = "findNamespace";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findNamespace_namespace_pathParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findNamespace_nsDescParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findNamespace_namespace_pathParamInfo {
            name            = "namespace_path";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findNamespace_nsDescParamInfo {
            name            = "nsDesc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sNamespaceInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTECSInfo_findRegionFunctionInfo {
            name            = "findRegion";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findRegion_namespace_pathParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findRegion_regionDescParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findRegion_namespace_pathParamInfo {
            name            = "namespace_path";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findRegion_regionDescParamInfo {
            name            = "regionDesc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sRegionInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTECSInfo_findSignatureFunctionInfo {
            name            = "findSignature";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findSignature_namespace_pathParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findSignature_signatureDescParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findSignature_namespace_pathParamInfo {
            name            = "namespace_path";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findSignature_signatureDescParamInfo {
            name            = "signatureDesc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sSignatureInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTECSInfo_findCelltypeFunctionInfo {
            name            = "findCelltype";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findCelltype_namespace_pathParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findCelltype_celltypeDescParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findCelltype_namespace_pathParamInfo {
            name            = "namespace_path";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findCelltype_celltypeDescParamInfo {
            name            = "celltypeDesc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sCelltypeInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTECSInfo_findCellFunctionInfo {
            name            = "findCell";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findCell_namespace_pathParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findCell_cellDescParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findCell_namespace_pathParamInfo {
            name            = "namespace_path";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findCell_cellDescParamInfo {
            name            = "cellDesc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sCellInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTECSInfo_findRawEntryDescriptorFunctionInfo {
            name            = "findRawEntryDescriptor";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findRawEntryDescriptor_namespace_pathParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findRawEntryDescriptor_rawEntryDescDescParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findRawEntryDescriptor_entryDescParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findRawEntryDescriptor_namespace_pathParamInfo {
            name            = "namespace_path";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findRawEntryDescriptor_rawEntryDescDescParamInfo {
            name            = "rawEntryDescDesc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sRawEntryDescriptorInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findRawEntryDescriptor_entryDescParamInfo {
            name            = "entryDesc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = Descriptor_of_nTECSInfo_sEntryInfo_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sTECSInfo_findRawEntryDescriptor_unsafeFunctionInfo {
            name            = "findRawEntryDescriptor_unsafe";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findRawEntryDescriptor_unsafe_namespace_pathParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findRawEntryDescriptor_unsafe_subscParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sTECSInfo_findRawEntryDescriptor_unsafe_rawDescParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findRawEntryDescriptor_unsafe_namespace_pathParamInfo {
            name            = "namespace_path";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findRawEntryDescriptor_unsafe_subscParamInfo {
            name            = "subsc";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sTECSInfo_findRawEntryDescriptor_unsafe_rawDescParamInfo {
            name            = "rawDesc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = void_Ptr__Ptr_TypeInfo.eTypeInfo;
        };

        /*** nTECSInfo_sAccessor signature information ****/
        cell nTECSInfo::tSignatureInfo nTECSInfo_sAccessorSignatureInfo {
            name            = "sAccessor";
            cFunctionInfo[] = nTECSInfo_sAccessor_selectNamespaceInfoByNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectCelltypeInfoByNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectSignatureInfoByNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectRegionInfoByNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectCellInfoByNameFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSignatureNameOfCellEntryFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedNamespaceInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectCelltypeInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectSignatureInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectNamespaceInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedCelltypeInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectCallInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectEntryInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectAttrInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectVarInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedAttrInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSizeIsExprOfAttrFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectTypeInfoOfAttrFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedVarInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSizeIsExprOfVarFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectTypeInfoOfVarFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedCallInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectSignatureOfCallFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedCallSpecifierInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedCallInternalInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedCallLocationInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedCallOptimizeInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedEntryInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectSignatureOfEntryFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedEntryInlineInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedSignatureInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectFunctionInfoByIndexFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedFunctionInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectTypeInfoOfReturnFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedParamInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectParamInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectTypeInfoOfParamFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedTypeInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectTypeInfoOfTypeFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedRegionInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectCellInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectRegionInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getSelectedCellInfoFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_selectCelltypeInfoOfCellFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getAttrValueInStrFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getAttrSizeIsValueFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getVarValueInStrFunctionInfo.eFunctionInfo;
            cFunctionInfo[] = nTECSInfo_sAccessor_getVarSizeIsValueFunctionInfo.eFunctionInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectNamespaceInfoByNameFunctionInfo {
            name            = "selectNamespaceInfoByName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectNamespaceInfoByName_namespacePathParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectNamespaceInfoByName_namespacePathParamInfo {
            name            = "namespacePath";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectCelltypeInfoByNameFunctionInfo {
            name            = "selectCelltypeInfoByName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectCelltypeInfoByName_celltypePathParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectCelltypeInfoByName_celltypePathParamInfo {
            name            = "celltypePath";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectSignatureInfoByNameFunctionInfo {
            name            = "selectSignatureInfoByName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectSignatureInfoByName_signaturePathParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectSignatureInfoByName_signaturePathParamInfo {
            name            = "signaturePath";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectRegionInfoByNameFunctionInfo {
            name            = "selectRegionInfoByName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectRegionInfoByName_regionPathParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectRegionInfoByName_regionPathParamInfo {
            name            = "regionPath";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectCellInfoByNameFunctionInfo {
            name            = "selectCellInfoByName";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectCellInfoByName_cellPathParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectCellInfoByName_cellPathParamInfo {
            name            = "cellPath";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSignatureNameOfCellEntryFunctionInfo {
            name            = "getSignatureNameOfCellEntry";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSignatureNameOfCellEntry_cellEntryPathParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSignatureNameOfCellEntry_signatureGlobalNameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSignatureNameOfCellEntry_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSignatureNameOfCellEntry_cellEntryPathParamInfo {
            name            = "cellEntryPath";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = "";
            cTypeInfo       = const__char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSignatureNameOfCellEntry_signatureGlobalNameParamInfo {
            name            = "signatureGlobalName";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $2";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSignatureNameOfCellEntry_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedNamespaceInfoFunctionInfo {
            name            = "getSelectedNamespaceInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedNamespaceInfo_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedNamespaceInfo_max_lenParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedNamespaceInfo_num_namespaceParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedNamespaceInfo_num_celltypeParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedNamespaceInfo_num_signatureParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedNamespaceInfo_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedNamespaceInfo_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedNamespaceInfo_num_namespaceParamInfo {
            name            = "num_namespace";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedNamespaceInfo_num_celltypeParamInfo {
            name            = "num_celltype";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedNamespaceInfo_num_signatureParamInfo {
            name            = "num_signature";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectCelltypeInfoFunctionInfo {
            name            = "selectCelltypeInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectCelltypeInfo_ithParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectCelltypeInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectSignatureInfoFunctionInfo {
            name            = "selectSignatureInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectSignatureInfo_ithParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectSignatureInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectNamespaceInfoFunctionInfo {
            name            = "selectNamespaceInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectNamespaceInfo_ithParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectNamespaceInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedCelltypeInfoFunctionInfo {
            name            = "getSelectedCelltypeInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCelltypeInfo_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCelltypeInfo_max_lenParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCelltypeInfo_num_attrParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCelltypeInfo_num_varParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCelltypeInfo_num_callParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCelltypeInfo_num_entryParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCelltypeInfo_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCelltypeInfo_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCelltypeInfo_num_attrParamInfo {
            name            = "num_attr";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCelltypeInfo_num_varParamInfo {
            name            = "num_var";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCelltypeInfo_num_callParamInfo {
            name            = "num_call";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCelltypeInfo_num_entryParamInfo {
            name            = "num_entry";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectCallInfoFunctionInfo {
            name            = "selectCallInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectCallInfo_ithParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectCallInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectEntryInfoFunctionInfo {
            name            = "selectEntryInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectEntryInfo_ithParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectEntryInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectAttrInfoFunctionInfo {
            name            = "selectAttrInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectAttrInfo_ithParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectAttrInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectVarInfoFunctionInfo {
            name            = "selectVarInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectVarInfo_ithParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectVarInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedAttrInfoFunctionInfo {
            name            = "getSelectedAttrInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedAttrInfo_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedAttrInfo_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedAttrInfo_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedAttrInfo_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSizeIsExprOfAttrFunctionInfo {
            name            = "getSizeIsExprOfAttr";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSizeIsExprOfAttr_expr_strParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSizeIsExprOfAttr_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSizeIsExprOfAttr_expr_strParamInfo {
            name            = "expr_str";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSizeIsExprOfAttr_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectTypeInfoOfAttrFunctionInfo {
            name            = "selectTypeInfoOfAttr";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedVarInfoFunctionInfo {
            name            = "getSelectedVarInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedVarInfo_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedVarInfo_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedVarInfo_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedVarInfo_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSizeIsExprOfVarFunctionInfo {
            name            = "getSizeIsExprOfVar";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSizeIsExprOfVar_expr_strParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSizeIsExprOfVar_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSizeIsExprOfVar_expr_strParamInfo {
            name            = "expr_str";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSizeIsExprOfVar_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectTypeInfoOfVarFunctionInfo {
            name            = "selectTypeInfoOfVar";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedCallInfoFunctionInfo {
            name            = "getSelectedCallInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallInfo_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallInfo_max_lenParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallInfo_array_sizeParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallInfo_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallInfo_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallInfo_array_sizeParamInfo {
            name            = "array_size";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectSignatureOfCallFunctionInfo {
            name            = "selectSignatureOfCall";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedCallSpecifierInfoFunctionInfo {
            name            = "getSelectedCallSpecifierInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallSpecifierInfo_b_optionalParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallSpecifierInfo_b_dynamicParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallSpecifierInfo_b_ref_descParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallSpecifierInfo_b_omitParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallSpecifierInfo_b_optionalParamInfo {
            name            = "b_optional";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallSpecifierInfo_b_dynamicParamInfo {
            name            = "b_dynamic";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallSpecifierInfo_b_ref_descParamInfo {
            name            = "b_ref_desc";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallSpecifierInfo_b_omitParamInfo {
            name            = "b_omit";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedCallInternalInfoFunctionInfo {
            name            = "getSelectedCallInternalInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallInternalInfo_b_allocator_portParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallInternalInfo_b_require_portParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallInternalInfo_b_allocator_portParamInfo {
            name            = "b_allocator_port";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallInternalInfo_b_require_portParamInfo {
            name            = "b_require_port";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedCallLocationInfoFunctionInfo {
            name            = "getSelectedCallLocationInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallLocationInfo_offsetParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallLocationInfo_placeParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallLocationInfo_offsetParamInfo {
            name            = "offset";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = uint32_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallLocationInfo_placeParamInfo {
            name            = "place";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int8_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedCallOptimizeInfoFunctionInfo {
            name            = "getSelectedCallOptimizeInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallOptimizeInfo_b_VMT_uselessParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallOptimizeInfo_b_skelton_uselessParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCallOptimizeInfo_b_cell_uniqueParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallOptimizeInfo_b_VMT_uselessParamInfo {
            name            = "b_VMT_useless";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallOptimizeInfo_b_skelton_uselessParamInfo {
            name            = "b_skelton_useless";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCallOptimizeInfo_b_cell_uniqueParamInfo {
            name            = "b_cell_unique";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedEntryInfoFunctionInfo {
            name            = "getSelectedEntryInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedEntryInfo_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedEntryInfo_max_lenParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedEntryInfo_array_sizeParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedEntryInfo_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedEntryInfo_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedEntryInfo_array_sizeParamInfo {
            name            = "array_size";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectSignatureOfEntryFunctionInfo {
            name            = "selectSignatureOfEntry";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedEntryInlineInfoFunctionInfo {
            name            = "getSelectedEntryInlineInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedEntryInlineInfo_b_inlineParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedEntryInlineInfo_b_inlineParamInfo {
            name            = "b_inline";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = bool_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedSignatureInfoFunctionInfo {
            name            = "getSelectedSignatureInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedSignatureInfo_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedSignatureInfo_max_lenParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedSignatureInfo_num_functionParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedSignatureInfo_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedSignatureInfo_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedSignatureInfo_num_functionParamInfo {
            name            = "num_function";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectFunctionInfoByIndexFunctionInfo {
            name            = "selectFunctionInfoByIndex";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectFunctionInfoByIndex_ithParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectFunctionInfoByIndex_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedFunctionInfoFunctionInfo {
            name            = "getSelectedFunctionInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedFunctionInfo_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedFunctionInfo_max_lenParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedFunctionInfo_num_argsParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedFunctionInfo_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedFunctionInfo_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedFunctionInfo_num_argsParamInfo {
            name            = "num_args";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectTypeInfoOfReturnFunctionInfo {
            name            = "selectTypeInfoOfReturn";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedParamInfoFunctionInfo {
            name            = "getSelectedParamInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedParamInfo_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedParamInfo_max_lenParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedParamInfo_dirParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedParamInfo_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedParamInfo_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedParamInfo_dirParamInfo {
            name            = "dir";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int8_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectParamInfoFunctionInfo {
            name            = "selectParamInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectParamInfo_ithParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectParamInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectTypeInfoOfParamFunctionInfo {
            name            = "selectTypeInfoOfParam";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedTypeInfoFunctionInfo {
            name            = "getSelectedTypeInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedTypeInfo_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedTypeInfo_max_lenParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedTypeInfo_kindParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedTypeInfo_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedTypeInfo_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedTypeInfo_kindParamInfo {
            name            = "kind";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int8_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectTypeInfoOfTypeFunctionInfo {
            name            = "selectTypeInfoOfType";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedRegionInfoFunctionInfo {
            name            = "getSelectedRegionInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedRegionInfo_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedRegionInfo_max_lenParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedRegionInfo_num_cellParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedRegionInfo_num_regionParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedRegionInfo_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedRegionInfo_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedRegionInfo_num_cellParamInfo {
            name            = "num_cell";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedRegionInfo_num_regionParamInfo {
            name            = "num_region";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectCellInfoFunctionInfo {
            name            = "selectCellInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectCellInfo_ithParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectCellInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectRegionInfoFunctionInfo {
            name            = "selectRegionInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_selectRegionInfo_ithParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_selectRegionInfo_ithParamInfo {
            name            = "ith";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getSelectedCellInfoFunctionInfo {
            name            = "getSelectedCellInfo";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCellInfo_nameParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getSelectedCellInfo_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCellInfo_nameParamInfo {
            name            = "name";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getSelectedCellInfo_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_selectCelltypeInfoOfCellFunctionInfo {
            name            = "selectCelltypeInfoOfCell";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getAttrValueInStrFunctionInfo {
            name            = "getAttrValueInStr";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getAttrValueInStr_bufParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getAttrValueInStr_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getAttrValueInStr_bufParamInfo {
            name            = "buf";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getAttrValueInStr_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getAttrSizeIsValueFunctionInfo {
            name            = "getAttrSizeIsValue";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getVarValueInStrFunctionInfo {
            name            = "getVarValueInStr";
            bOneway         = false;
            cParamInfo[]    = nTECSInfo_sAccessor_getVarValueInStr_bufParamInfo.eParamInfo;
            cParamInfo[]    = nTECSInfo_sAccessor_getVarValueInStr_max_lenParamInfo.eParamInfo;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getVarValueInStr_bufParamInfo {
            name            = "buf";
            dir             = PARAM_DIR_OUT;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = " $1";
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tParamInfo nTECSInfo_sAccessor_getVarValueInStr_max_lenParamInfo {
            name            = "max_len";
            dir             = PARAM_DIR_IN;
            sizeIsExpr      = (char_t*)0;
            countIsExpr     = (char_t*)0;
            stringExpr      = (char_t*)0;
            cTypeInfo       = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tFunctionInfo nTECSInfo_sAccessor_getVarSizeIsValueFunctionInfo {
            name            = "getVarSizeIsValue";
            bOneway         = false;
            cReturnTypeInfo = ERTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tCelltypeInfo nTECSInfo_tTECSInfoCelltypeInfo {
            name             = "tTECSInfo";
            b_singleton      = true;
            b_IDX_is_ID_act  = C_EXP( "nTECSInfo_tTECSInfo__IDX_is_ID_act" );
            sizeOfCB         = C_EXP( "nTECSInfo_tTECSInfo__sizeOfCB" );
            sizeOfINIB       = C_EXP( "nTECSInfo_tTECSInfo__sizeOfINIB" );
            n_cellInLinkUnit = C_EXP( "nTECSInfo_tTECSInfo__NCELLINLINKUNIT" );
            n_cellInSystem   = 1;
            cEntryInfo[]    = nTECSInfo_tTECSInfo_eTECSInfoEntryInfo.eEntryInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfo_cTECSInfoCallInfo.eCallInfo;
        };
        cell nTECSInfo::tEntryInfo nTECSInfo_tTECSInfo_eTECSInfoEntryInfo{
            name            = "eTECSInfo";
            cSignatureInfo  = nTECSInfo_sTECSInfoSignatureInfo.eSignatureInfo;
            b_inline        = true;
            array_size      = C_EXP( "nTECSInfo_tTECSInfo_eTECSInfo__array_size" );
        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfo_cTECSInfoCallInfo{
            name            = "cTECSInfo";
            cSignatureInfo  = nTECSInfo_sTECSInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfo_cTECSInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfo_cTECSInfo__array_size" );
            b_optional        = false;
            b_omit            = false;
            b_dynamic         = false;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfo_cTECSInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfo_cTECSInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfo_cTECSInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfo_cTECSInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCelltypeInfo nTECSInfo_tTECSInfoAccessorCelltypeInfo {
            name             = "tTECSInfoAccessor";
            b_singleton      = false;
            b_IDX_is_ID_act  = C_EXP( "nTECSInfo_tTECSInfoAccessor__IDX_is_ID_act" );
            sizeOfCB         = C_EXP( "nTECSInfo_tTECSInfoAccessor__sizeOfCB" );
            sizeOfINIB       = C_EXP( "nTECSInfo_tTECSInfoAccessor__sizeOfINIB" );
            n_cellInLinkUnit = C_EXP( "nTECSInfo_tTECSInfoAccessor__NCELLINLINKUNIT" );
            n_cellInSystem   = 1;
            cEntryInfo[]    = nTECSInfo_tTECSInfoAccessor_eSelectorEntryInfo.eEntryInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cTECSInfoCallInfo.eCallInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cNSInfoCallInfo.eCallInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cCelltypeInfoCallInfo.eCallInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cSignatureInfoCallInfo.eCallInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cFunctionInfoCallInfo.eCallInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cParamInfoCallInfo.eCallInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cCallInfoCallInfo.eCallInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cEntryInfoCallInfo.eCallInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cAttrInfoCallInfo.eCallInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cVarInfoCallInfo.eCallInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cVarDeclInfoCallInfo.eCallInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cTypeInfoCallInfo.eCallInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cRegionInfoCallInfo.eCallInfo;
            cCallInfo[]     = nTECSInfo_tTECSInfoAccessor_cCellInfoCallInfo.eCallInfo;
            cAttrInfo[]     = nTECSInfo_tTECSInfoAccessor_NAME_LENVarDeclInfo.eVarDeclInfo;
            cVarInfo[]      = nTECSInfo_tTECSInfoAccessor_nameVarDeclInfo.eVarDeclInfo;
            cVarInfo[]      = nTECSInfo_tTECSInfoAccessor_name2VarDeclInfo.eVarDeclInfo;
            cVarInfo[]      = nTECSInfo_tTECSInfoAccessor_selectedCbpVarDeclInfo.eVarDeclInfo;
            cVarInfo[]      = nTECSInfo_tTECSInfoAccessor_selectedInibpVarDeclInfo.eVarDeclInfo;
            cVarInfo[]      = nTECSInfo_tTECSInfoAccessor_TDescVarDeclInfo.eVarDeclInfo;
        };
        cell nTECSInfo::tEntryInfo nTECSInfo_tTECSInfoAccessor_eSelectorEntryInfo{
            name            = "eSelector";
            cSignatureInfo  = nTECSInfo_sAccessorSignatureInfo.eSignatureInfo;
            b_inline        = false;
            array_size      = C_EXP( "nTECSInfo_tTECSInfoAccessor_eSelector__array_size" );
        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cTECSInfoCallInfo{
            name            = "cTECSInfo";
            cSignatureInfo  = nTECSInfo_sTECSInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cTECSInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cTECSInfo__array_size" );
            b_optional        = false;
            b_omit            = false;
            b_dynamic         = false;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cTECSInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cTECSInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cTECSInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cTECSInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cNSInfoCallInfo{
            name            = "cNSInfo";
            cSignatureInfo  = nTECSInfo_sNamespaceInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cNSInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cNSInfo__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = true;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cNSInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cNSInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cNSInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cNSInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cCelltypeInfoCallInfo{
            name            = "cCelltypeInfo";
            cSignatureInfo  = nTECSInfo_sCelltypeInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCelltypeInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCelltypeInfo__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = true;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCelltypeInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCelltypeInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCelltypeInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCelltypeInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cSignatureInfoCallInfo{
            name            = "cSignatureInfo";
            cSignatureInfo  = nTECSInfo_sSignatureInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cSignatureInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cSignatureInfo__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = true;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cSignatureInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cSignatureInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cSignatureInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cSignatureInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cFunctionInfoCallInfo{
            name            = "cFunctionInfo";
            cSignatureInfo  = nTECSInfo_sFunctionInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cFunctionInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cFunctionInfo__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = true;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cFunctionInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cFunctionInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cFunctionInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cFunctionInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cParamInfoCallInfo{
            name            = "cParamInfo";
            cSignatureInfo  = nTECSInfo_sParamInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cParamInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cParamInfo__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = true;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cParamInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cParamInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cParamInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cParamInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cCallInfoCallInfo{
            name            = "cCallInfo";
            cSignatureInfo  = nTECSInfo_sCallInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCallInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCallInfo__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = true;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCallInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCallInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCallInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCallInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cEntryInfoCallInfo{
            name            = "cEntryInfo";
            cSignatureInfo  = nTECSInfo_sEntryInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cEntryInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cEntryInfo__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = true;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cEntryInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cEntryInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cEntryInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cEntryInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cAttrInfoCallInfo{
            name            = "cAttrInfo";
            cSignatureInfo  = nTECSInfo_sVarDeclInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cAttrInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cAttrInfo__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = true;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cAttrInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cAttrInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cAttrInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cAttrInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cVarInfoCallInfo{
            name            = "cVarInfo";
            cSignatureInfo  = nTECSInfo_sVarDeclInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cVarInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cVarInfo__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = true;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cVarInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cVarInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cVarInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cVarInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cVarDeclInfoCallInfo{
            name            = "cVarDeclInfo";
            cSignatureInfo  = nTECSInfo_sVarDeclInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cVarDeclInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cVarDeclInfo__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = true;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cVarDeclInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cVarDeclInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cVarDeclInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cVarDeclInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cTypeInfoCallInfo{
            name            = "cTypeInfo";
            cSignatureInfo  = nTECSInfo_sTypeInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cTypeInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cTypeInfo__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = true;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cTypeInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cTypeInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cTypeInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cTypeInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cRegionInfoCallInfo{
            name            = "cRegionInfo";
            cSignatureInfo  = nTECSInfo_sRegionInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cRegionInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cRegionInfo__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = true;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cRegionInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cRegionInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cRegionInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cRegionInfo__b_cell_unique" );

        };
        cell nTECSInfo::tCallInfo nTECSInfo_tTECSInfoAccessor_cCellInfoCallInfo{
            name            = "cCellInfo";
            cSignatureInfo  = nTECSInfo_sCellInfoSignatureInfo.eSignatureInfo;
            offset            = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCellInfo__offset" );
            array_size        = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCellInfo__array_size" );
            b_optional        = true;
            b_omit            = false;
            b_dynamic         = true;
            b_ref_desc        = false;
            b_allocator_port  = false;
            b_require_port    = false;
            place             = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCellInfo__place" );
            b_VMT_useless     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCellInfo__b_VMT_useless" );
            b_skelton_useless = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCellInfo__b_skelton_useless" );
            b_cell_unique     = C_EXP( "nTECSInfo_tTECSInfoAccessor_cCellInfo__b_cell_unique" );

        };
        cell nTECSInfo::tVarDeclInfo nTECSInfo_tTECSInfoAccessor_NAME_LENVarDeclInfo {
            name            = "NAME_LEN";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_ATTR;
            offset          = C_EXP( "OFFSET_OF_nTECSInfo_tTECSInfoAccessor_NAME_LEN" );
            place           = C_EXP( "PLACE_OF_nTECSInfo_tTECSInfoAccessor_NAME_LEN" );
            cTypeInfo       = int16_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo nTECSInfo_tTECSInfoAccessor_nameVarDeclInfo {
            name            = "name";
            sizeIsExpr      = "mikan";
            declType        = DECLTYPE_VAR;
            offset          = C_EXP( "OFFSET_OF_nTECSInfo_tTECSInfoAccessor_name" );
            place           = C_EXP( "PLACE_OF_nTECSInfo_tTECSInfoAccessor_name" );
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo nTECSInfo_tTECSInfoAccessor_name2VarDeclInfo {
            name            = "name2";
            sizeIsExpr      = "mikan";
            declType        = DECLTYPE_VAR;
            offset          = C_EXP( "OFFSET_OF_nTECSInfo_tTECSInfoAccessor_name2" );
            place           = C_EXP( "PLACE_OF_nTECSInfo_tTECSInfoAccessor_name2" );
            cTypeInfo       = char_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo nTECSInfo_tTECSInfoAccessor_selectedCbpVarDeclInfo {
            name            = "selectedCbp";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_VAR;
            offset          = C_EXP( "OFFSET_OF_nTECSInfo_tTECSInfoAccessor_selectedCbp" );
            place           = C_EXP( "PLACE_OF_nTECSInfo_tTECSInfoAccessor_selectedCbp" );
            cTypeInfo       = int8_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo nTECSInfo_tTECSInfoAccessor_selectedInibpVarDeclInfo {
            name            = "selectedInibp";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_VAR;
            offset          = C_EXP( "OFFSET_OF_nTECSInfo_tTECSInfoAccessor_selectedInibp" );
            place           = C_EXP( "PLACE_OF_nTECSInfo_tTECSInfoAccessor_selectedInibp" );
            cTypeInfo       = int8_t_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVarDeclInfo nTECSInfo_tTECSInfoAccessor_TDescVarDeclInfo {
            name            = "TDesc";
            sizeIsExpr      = (char_t*)0;
            declType        = DECLTYPE_VAR;
            offset          = C_EXP( "OFFSET_OF_nTECSInfo_tTECSInfoAccessor_TDesc" );
            place           = C_EXP( "PLACE_OF_nTECSInfo_tTECSInfoAccessor_TDesc" );
            cTypeInfo       = Descriptor_of_nTECSInfo_sTypeInfoTypeInfo.eTypeInfo;
        };

        /*** :: region information cell ***/
        cell nTECSInfo::tRegionInfo _LinkRootRegionInfo{
            name = "::";
            cCellInfo[] = PutStringStdioCellInfo.eCellInfo;
            cCellInfo[] = HelloWorldCellInfo.eCellInfo;
            cRegionInfo[] = rTEMPRegionInfo.eRegionInfo;
        };

        /*** PutStringStdio cell information ****/
        cell nTECSInfo::tCellInfo PutStringStdioCellInfo {
            name            = "PutStringStdio";
            cbp             = C_EXP( "PutStringStdio__CBP" );
            inibp           = C_EXP( "PutStringStdio__INIBP" );
            cCelltypeInfo   = tPutStringStdioCelltypeInfo.eCelltypeInfo;
            cRawEntryDescriptor[] = PutStringStdio_ePutStringRawEntryDescriptorInfo.eRawEntryDescriptor;
        };
        cell nTECSInfo::tRawEntryDescriptorInfo PutStringStdio_ePutStringRawEntryDescriptorInfo {
           size = 1;
           rawEntryDescriptor = { C_EXP( "&PutStringStdio_ePutString_des" ) };
        };

        /*** HelloWorld cell information ****/
        cell nTECSInfo::tCellInfo HelloWorldCellInfo {
            name            = "HelloWorld";
            cbp             = C_EXP( "HelloWorld__CBP" );
            inibp           = C_EXP( "HelloWorld__INIBP" );
            cCelltypeInfo   = tHelloWorldCelltypeInfo.eCelltypeInfo;
            cRawEntryDescriptor[] = HelloWorld_eMainRawEntryDescriptorInfo.eRawEntryDescriptor;
        };
        cell nTECSInfo::tRawEntryDescriptorInfo HelloWorld_eMainRawEntryDescriptorInfo {
           size = 1;
           rawEntryDescriptor = { C_EXP( "&HelloWorld_eMain_des" ) };
        };

        /*** ::rTEMP region information cell ***/
        cell nTECSInfo::tRegionInfo rTEMPRegionInfo{
            name = "rTEMP";
            cCellInfo[] = rTEMP_TaskCellInfo.eCellInfo;
            cCellInfo[] = rTEMP_TaskMainCellInfo.eCellInfo;
            cCellInfo[] = rTEMP_TECSInfoCompo_TECSInfoCellInfo.eCellInfo;
            cCellInfo[] = rTEMP_TECSInfoCompo_TECSInfoAccessorCellInfo.eCellInfo;
            cRegionInfo[] = rTEMP_rTECSInfoRegionInfo.eRegionInfo;
        };

        /*** rTEMP_Task cell information ****/
        cell nTECSInfo::tCellInfo rTEMP_TaskCellInfo {
            name            = "Task";
            cbp             = C_EXP( "rTEMP_Task__CBP" );
            inibp           = C_EXP( "rTEMP_Task__INIBP" );
            cCelltypeInfo   = tTaskCelltypeInfo.eCelltypeInfo;
            cRawEntryDescriptor[] = rTEMP_Task_eTaskRawEntryDescriptorInfo.eRawEntryDescriptor;
        };
        cell nTECSInfo::tRawEntryDescriptorInfo rTEMP_Task_eTaskRawEntryDescriptorInfo {
           size = 1;
           rawEntryDescriptor = { C_EXP( "&rTEMP_Task_eTask_des" ) };
        };

        /*** rTEMP_TaskMain cell information ****/
        cell nTECSInfo::tCellInfo rTEMP_TaskMainCellInfo {
            name            = "TaskMain";
            cbp             = C_EXP( "rTEMP_TaskMain__CBP" );
            inibp           = C_EXP( "rTEMP_TaskMain__INIBP" );
            cCelltypeInfo   = tTaskMainCelltypeInfo.eCelltypeInfo;
            cRawEntryDescriptor[] = rTEMP_TaskMain_eBodyRawEntryDescriptorInfo.eRawEntryDescriptor;
        };
        cell nTECSInfo::tRawEntryDescriptorInfo rTEMP_TaskMain_eBodyRawEntryDescriptorInfo {
           size = 1;
           rawEntryDescriptor = { C_EXP( "&rTEMP_TaskMain_eBody_des" ) };
        };

        /*** rTEMP_TECSInfoCompo_TECSInfo cell information ****/
        cell nTECSInfo::tCellInfo rTEMP_TECSInfoCompo_TECSInfoCellInfo {
            name            = "TECSInfoCompo_TECSInfo";
            cbp             = C_EXP( "rTEMP_TECSInfoCompo_TECSInfo__CBP" );
            inibp           = C_EXP( "rTEMP_TECSInfoCompo_TECSInfo__INIBP" );
            cCelltypeInfo   = nTECSInfo_tTECSInfoCelltypeInfo.eCelltypeInfo;
            cRawEntryDescriptor[] = rTEMP_TECSInfoCompo_TECSInfo_eTECSInfoRawEntryDescriptorInfo.eRawEntryDescriptor;
        };
        cell nTECSInfo::tRawEntryDescriptorInfo rTEMP_TECSInfoCompo_TECSInfo_eTECSInfoRawEntryDescriptorInfo {
           size = 1;
           rawEntryDescriptor = { C_EXP( "&rTEMP_TECSInfoCompo_TECSInfo_eTECSInfo_des" ) };
        };

        /*** rTEMP_TECSInfoCompo_TECSInfoAccessor cell information ****/
        cell nTECSInfo::tCellInfo rTEMP_TECSInfoCompo_TECSInfoAccessorCellInfo {
            name            = "TECSInfoCompo_TECSInfoAccessor";
            cbp             = C_EXP( "rTEMP_TECSInfoCompo_TECSInfoAccessor__CBP" );
            inibp           = C_EXP( "rTEMP_TECSInfoCompo_TECSInfoAccessor__INIBP" );
            cCelltypeInfo   = nTECSInfo_tTECSInfoAccessorCelltypeInfo.eCelltypeInfo;
            cRawEntryDescriptor[] = rTEMP_TECSInfoCompo_TECSInfoAccessor_eSelectorRawEntryDescriptorInfo.eRawEntryDescriptor;
        };
        cell nTECSInfo::tRawEntryDescriptorInfo rTEMP_TECSInfoCompo_TECSInfoAccessor_eSelectorRawEntryDescriptorInfo {
           size = 1;
           rawEntryDescriptor = { C_EXP( "&rTEMP_TECSInfoCompo_TECSInfoAccessor_eSelector_des" ) };
        };

        /*** ::rTEMP::rTECSInfo region information cell ***/
        cell nTECSInfo::tRegionInfo rTEMP_rTECSInfoRegionInfo{
            name = "rTECSInfo";
        };

        /*** TYPE information cell ***/
        cell nTECSInfo::tVoidTypeInfo voidTypeInfo{
            name           = "void";
            typeKind       = TECSTypeKind_VoidType;
            size           = C_EXP( "sizeof(void)" );
            b_const        = false;
            b_volatile     = false;
        };
        cell nTECSInfo::tDefinedTypeInfo TEXPTNTypeInfo{
            name           = "TEXPTN";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(TEXPTN)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = uint_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo uint_tTypeInfo{
            name           = "uint_t";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(uint_t)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = unsigned__intTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tIntTypeInfo unsigned__intTypeInfo{
            name           = "unsigned int";
            typeKind       = TECSTypeKind_IntType;
            size           = C_EXP( "sizeof(unsigned int)" );
            b_const        = false;
            b_volatile     = false;
        };
        cell nTECSInfo::tDefinedTypeInfo ERTypeInfo{
            name           = "ER";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(ER)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo int_tTypeInfo{
            name           = "int_t";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(int_t)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = signed__intTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tIntTypeInfo signed__intTypeInfo{
            name           = "signed int";
            typeKind       = TECSTypeKind_IntType;
            size           = C_EXP( "sizeof(signed int)" );
            b_const        = false;
            b_volatile     = false;
        };
        cell nTECSInfo::tDefinedTypeInfo RELTIMTypeInfo{
            name           = "RELTIM";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(RELTIM)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = uint_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tPtrTypeInfo SYSTIM_Ptr_TypeInfo{
            name           = "SYSTIM*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(SYSTIM*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = SYSTIMTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo SYSTIMTypeInfo{
            name           = "SYSTIM";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(SYSTIM)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = ulong_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo ulong_tTypeInfo{
            name           = "ulong_t";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(ulong_t)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = unsigned__longTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tIntTypeInfo unsigned__longTypeInfo{
            name           = "unsigned long";
            typeKind       = TECSTypeKind_IntType;
            size           = C_EXP( "sizeof(unsigned long)" );
            b_const        = false;
            b_volatile     = false;
        };
        cell nTECSInfo::tPtrTypeInfo SYSUTM_Ptr_TypeInfo{
            name           = "SYSUTM*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(SYSUTM*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = SYSUTMTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo SYSUTMTypeInfo{
            name           = "SYSUTM";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(SYSUTM)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = ulong_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo TMOTypeInfo{
            name           = "TMO";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(TMO)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tPtrTypeInfo T_RSEM_Ptr_TypeInfo{
            name           = "T_RSEM*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(T_RSEM*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = T_RSEMTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo T_RSEMTypeInfo{
            name           = "T_RSEM";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(T_RSEM)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = struct__t_rsemTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tStructTypeInfo struct__t_rsemTypeInfo{
            name           = "struct t_rsem";
            typeKind       = TECSTypeKind_StructType;
            size           = C_EXP( "sizeof(struct t_rsem)" );
            b_const        = false;
            b_volatile     = false;
            cVarDeclInfo[] = struct__t_rsem_wtskidVarDeclInfo.eVarDeclInfo;
            cVarDeclInfo[] = struct__t_rsem_semcntVarDeclInfo.eVarDeclInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo IDTypeInfo{
            name           = "ID";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(ID)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo FLGPTNTypeInfo{
            name           = "FLGPTN";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(FLGPTN)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = uint_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo MODETypeInfo{
            name           = "MODE";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(MODE)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = uint_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tPtrTypeInfo FLGPTN_Ptr_TypeInfo{
            name           = "FLGPTN*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(FLGPTN*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = FLGPTNTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tPtrTypeInfo T_RFLG_Ptr_TypeInfo{
            name           = "T_RFLG*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(T_RFLG*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = T_RFLGTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo T_RFLGTypeInfo{
            name           = "T_RFLG";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(T_RFLG)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = struct__t_rflgTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tStructTypeInfo struct__t_rflgTypeInfo{
            name           = "struct t_rflg";
            typeKind       = TECSTypeKind_StructType;
            size           = C_EXP( "sizeof(struct t_rflg)" );
            b_const        = false;
            b_volatile     = false;
            cVarDeclInfo[] = struct__t_rflg_wtskidVarDeclInfo.eVarDeclInfo;
            cVarDeclInfo[] = struct__t_rflg_flgptnVarDeclInfo.eVarDeclInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo intptr_tTypeInfo{
            name           = "intptr_t";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(intptr_t)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = longTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tIntTypeInfo longTypeInfo{
            name           = "long";
            typeKind       = TECSTypeKind_IntType;
            size           = C_EXP( "sizeof(long)" );
            b_const        = false;
            b_volatile     = false;
        };
        cell nTECSInfo::tPtrTypeInfo intptr_t_Ptr_TypeInfo{
            name           = "intptr_t*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(intptr_t*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = intptr_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tPtrTypeInfo T_RDTQ_Ptr_TypeInfo{
            name           = "T_RDTQ*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(T_RDTQ*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = T_RDTQTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo T_RDTQTypeInfo{
            name           = "T_RDTQ";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(T_RDTQ)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = struct__t_rdtqTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tStructTypeInfo struct__t_rdtqTypeInfo{
            name           = "struct t_rdtq";
            typeKind       = TECSTypeKind_StructType;
            size           = C_EXP( "sizeof(struct t_rdtq)" );
            b_const        = false;
            b_volatile     = false;
            cVarDeclInfo[] = struct__t_rdtq_stskidVarDeclInfo.eVarDeclInfo;
            cVarDeclInfo[] = struct__t_rdtq_rtskidVarDeclInfo.eVarDeclInfo;
            cVarDeclInfo[] = struct__t_rdtq_sdtqcntVarDeclInfo.eVarDeclInfo;
        };
        cell nTECSInfo::tPtrTypeInfo const__char_t_Ptr_TypeInfo{
            name           = "const char_t*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(const char_t*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = const__char_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tIntTypeInfo const__char_tTypeInfo{
            name           = "const char_t";
            typeKind       = TECSTypeKind_IntType;
            size           = C_EXP( "sizeof(const char_t)" );
            b_const        = true;
            b_volatile     = false;
        };
        cell nTECSInfo::tDefinedTypeInfo ATRTypeInfo{
            name           = "ATR";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(ATR)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = uint_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo PRITypeInfo{
            name           = "PRI";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(PRI)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = int_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo size_tTypeInfo{
            name           = "size_t";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(size_t)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = unsigned__longTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tPtrTypeInfo char_t_Ptr_TypeInfo{
            name           = "char_t*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(char_t*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = char_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tIntTypeInfo char_tTypeInfo{
            name           = "char_t";
            typeKind       = TECSTypeKind_IntType;
            size           = C_EXP( "sizeof(char_t)" );
            b_const        = false;
            b_volatile     = false;
        };
        cell nTECSInfo::tDefinedTypeInfo pthread_tTypeInfo{
            name           = "pthread_t";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(pthread_t)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = intptr_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo pthread_cond_tTypeInfo{
            name           = "pthread_cond_t";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(pthread_cond_t)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = intptr_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDefinedTypeInfo pthread_mutex_tTypeInfo{
            name           = "pthread_mutex_t";
            typeKind       = TECSTypeKind_DefinedType;
            size           = C_EXP( "sizeof(pthread_mutex_t)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = intptr_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tIntTypeInfo int16_tTypeInfo{
            name           = "int16_t";
            typeKind       = TECSTypeKind_IntType;
            size           = C_EXP( "sizeof(int16_t)" );
            b_const        = false;
            b_volatile     = false;
        };
        cell nTECSInfo::tIntTypeInfo uint16_tTypeInfo{
            name           = "uint16_t";
            typeKind       = TECSTypeKind_IntType;
            size           = C_EXP( "sizeof(uint16_t)" );
            b_const        = false;
            b_volatile     = false;
        };
        cell nTECSInfo::tIntTypeInfo uint32_tTypeInfo{
            name           = "uint32_t";
            typeKind       = TECSTypeKind_IntType;
            size           = C_EXP( "sizeof(uint32_t)" );
            b_const        = false;
            b_volatile     = false;
        };
        cell nTECSInfo::tIntTypeInfo int8_tTypeInfo{
            name           = "int8_t";
            typeKind       = TECSTypeKind_IntType;
            size           = C_EXP( "sizeof(int8_t)" );
            b_const        = false;
            b_volatile     = false;
        };
        cell nTECSInfo::tPtrTypeInfo Descriptor_of_nTECSInfo_sTypeInfo_Ptr_TypeInfo{
            name           = "Descriptor( nTECSInfo_sTypeInfo )*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sTypeInfo )*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = Descriptor_of_nTECSInfo_sTypeInfoTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDescriptorTypeInfo Descriptor_of_nTECSInfo_sTypeInfoTypeInfo{
            name           = "Descriptor( nTECSInfo_sTypeInfo )";
            typeKind       = TECSTypeKind_DescriptorType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sTypeInfo ))" );
            b_const        = false;
            b_volatile     = false;
            cSignatureInfo   = nTECSInfo_sTypeInfoSignatureInfo.eSignatureInfo;
        };
        cell nTECSInfo::tPtrTypeInfo Descriptor_of_nTECSInfo_sVarDeclInfo_Ptr_TypeInfo{
            name           = "Descriptor( nTECSInfo_sVarDeclInfo )*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sVarDeclInfo )*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = Descriptor_of_nTECSInfo_sVarDeclInfoTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDescriptorTypeInfo Descriptor_of_nTECSInfo_sVarDeclInfoTypeInfo{
            name           = "Descriptor( nTECSInfo_sVarDeclInfo )";
            typeKind       = TECSTypeKind_DescriptorType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sVarDeclInfo ))" );
            b_const        = false;
            b_volatile     = false;
            cSignatureInfo   = nTECSInfo_sVarDeclInfoSignatureInfo.eSignatureInfo;
        };
        cell nTECSInfo::tPtrTypeInfo uint32_t_Ptr_TypeInfo{
            name           = "uint32_t*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(uint32_t*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = uint32_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tPtrTypeInfo int8_t_Ptr_TypeInfo{
            name           = "int8_t*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(int8_t*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = int8_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tIntTypeInfo int32_tTypeInfo{
            name           = "int32_t";
            typeKind       = TECSTypeKind_IntType;
            size           = C_EXP( "sizeof(int32_t)" );
            b_const        = false;
            b_volatile     = false;
        };
        cell nTECSInfo::tPtrTypeInfo const__void_Ptr_TypeInfo{
            name           = "const void*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(const void*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = const__voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tVoidTypeInfo const__voidTypeInfo{
            name           = "const void";
            typeKind       = TECSTypeKind_VoidType;
            size           = C_EXP( "sizeof(const void)" );
            b_const        = true;
            b_volatile     = false;
        };
        cell nTECSInfo::tPtrTypeInfo Descriptor_of_nTECSInfo_sParamInfo_Ptr_TypeInfo{
            name           = "Descriptor( nTECSInfo_sParamInfo )*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sParamInfo )*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = Descriptor_of_nTECSInfo_sParamInfoTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDescriptorTypeInfo Descriptor_of_nTECSInfo_sParamInfoTypeInfo{
            name           = "Descriptor( nTECSInfo_sParamInfo )";
            typeKind       = TECSTypeKind_DescriptorType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sParamInfo ))" );
            b_const        = false;
            b_volatile     = false;
            cSignatureInfo   = nTECSInfo_sParamInfoSignatureInfo.eSignatureInfo;
        };
        cell nTECSInfo::tPtrTypeInfo Descriptor_of_nTECSInfo_sFunctionInfo_Ptr_TypeInfo{
            name           = "Descriptor( nTECSInfo_sFunctionInfo )*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sFunctionInfo )*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = Descriptor_of_nTECSInfo_sFunctionInfoTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDescriptorTypeInfo Descriptor_of_nTECSInfo_sFunctionInfoTypeInfo{
            name           = "Descriptor( nTECSInfo_sFunctionInfo )";
            typeKind       = TECSTypeKind_DescriptorType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sFunctionInfo ))" );
            b_const        = false;
            b_volatile     = false;
            cSignatureInfo   = nTECSInfo_sFunctionInfoSignatureInfo.eSignatureInfo;
        };
        cell nTECSInfo::tPtrTypeInfo Descriptor_of_nTECSInfo_sSignatureInfo_Ptr_TypeInfo{
            name           = "Descriptor( nTECSInfo_sSignatureInfo )*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sSignatureInfo )*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = Descriptor_of_nTECSInfo_sSignatureInfoTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDescriptorTypeInfo Descriptor_of_nTECSInfo_sSignatureInfoTypeInfo{
            name           = "Descriptor( nTECSInfo_sSignatureInfo )";
            typeKind       = TECSTypeKind_DescriptorType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sSignatureInfo ))" );
            b_const        = false;
            b_volatile     = false;
            cSignatureInfo   = nTECSInfo_sSignatureInfoSignatureInfo.eSignatureInfo;
        };
        cell nTECSInfo::tPtrTypeInfo bool_t_Ptr_TypeInfo{
            name           = "bool_t*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(bool_t*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = bool_tTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tBoolTypeInfo bool_tTypeInfo{
            name           = "bool_t";
            typeKind       = TECSTypeKind_BoolType;
            size           = C_EXP( "sizeof(bool_t)" );
            b_const        = false;
            b_volatile     = false;
        };
        cell nTECSInfo::tPtrTypeInfo Descriptor_of_nTECSInfo_sCallInfo_Ptr_TypeInfo{
            name           = "Descriptor( nTECSInfo_sCallInfo )*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sCallInfo )*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = Descriptor_of_nTECSInfo_sCallInfoTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDescriptorTypeInfo Descriptor_of_nTECSInfo_sCallInfoTypeInfo{
            name           = "Descriptor( nTECSInfo_sCallInfo )";
            typeKind       = TECSTypeKind_DescriptorType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sCallInfo ))" );
            b_const        = false;
            b_volatile     = false;
            cSignatureInfo   = nTECSInfo_sCallInfoSignatureInfo.eSignatureInfo;
        };
        cell nTECSInfo::tPtrTypeInfo Descriptor_of_nTECSInfo_sEntryInfo_Ptr_TypeInfo{
            name           = "Descriptor( nTECSInfo_sEntryInfo )*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sEntryInfo )*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = Descriptor_of_nTECSInfo_sEntryInfoTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDescriptorTypeInfo Descriptor_of_nTECSInfo_sEntryInfoTypeInfo{
            name           = "Descriptor( nTECSInfo_sEntryInfo )";
            typeKind       = TECSTypeKind_DescriptorType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sEntryInfo ))" );
            b_const        = false;
            b_volatile     = false;
            cSignatureInfo   = nTECSInfo_sEntryInfoSignatureInfo.eSignatureInfo;
        };
        cell nTECSInfo::tPtrTypeInfo Descriptor_of_nTECSInfo_sRawEntryDescriptorInfo_Ptr_TypeInfo{
            name           = "Descriptor( nTECSInfo_sRawEntryDescriptorInfo )*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sRawEntryDescriptorInfo )*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = Descriptor_of_nTECSInfo_sRawEntryDescriptorInfoTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDescriptorTypeInfo Descriptor_of_nTECSInfo_sRawEntryDescriptorInfoTypeInfo{
            name           = "Descriptor( nTECSInfo_sRawEntryDescriptorInfo )";
            typeKind       = TECSTypeKind_DescriptorType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sRawEntryDescriptorInfo ))" );
            b_const        = false;
            b_volatile     = false;
            cSignatureInfo   = nTECSInfo_sRawEntryDescriptorInfoSignatureInfo.eSignatureInfo;
        };
        cell nTECSInfo::tPtrTypeInfo Descriptor_of_nTECSInfo_sCelltypeInfo_Ptr_TypeInfo{
            name           = "Descriptor( nTECSInfo_sCelltypeInfo )*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sCelltypeInfo )*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = Descriptor_of_nTECSInfo_sCelltypeInfoTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDescriptorTypeInfo Descriptor_of_nTECSInfo_sCelltypeInfoTypeInfo{
            name           = "Descriptor( nTECSInfo_sCelltypeInfo )";
            typeKind       = TECSTypeKind_DescriptorType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sCelltypeInfo ))" );
            b_const        = false;
            b_volatile     = false;
            cSignatureInfo   = nTECSInfo_sCelltypeInfoSignatureInfo.eSignatureInfo;
        };
        cell nTECSInfo::tPtrTypeInfo void_Ptr__Ptr_TypeInfo{
            name           = "void**";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(void**)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = void_Ptr_TypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tPtrTypeInfo void_Ptr_TypeInfo{
            name           = "void*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(void*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = voidTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tPtrTypeInfo Descriptor_of_nTECSInfo_sNamespaceInfo_Ptr_TypeInfo{
            name           = "Descriptor( nTECSInfo_sNamespaceInfo )*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sNamespaceInfo )*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = Descriptor_of_nTECSInfo_sNamespaceInfoTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDescriptorTypeInfo Descriptor_of_nTECSInfo_sNamespaceInfoTypeInfo{
            name           = "Descriptor( nTECSInfo_sNamespaceInfo )";
            typeKind       = TECSTypeKind_DescriptorType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sNamespaceInfo ))" );
            b_const        = false;
            b_volatile     = false;
            cSignatureInfo   = nTECSInfo_sNamespaceInfoSignatureInfo.eSignatureInfo;
        };
        cell nTECSInfo::tPtrTypeInfo Descriptor_of_nTECSInfo_sCellInfo_Ptr_TypeInfo{
            name           = "Descriptor( nTECSInfo_sCellInfo )*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sCellInfo )*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = Descriptor_of_nTECSInfo_sCellInfoTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDescriptorTypeInfo Descriptor_of_nTECSInfo_sCellInfoTypeInfo{
            name           = "Descriptor( nTECSInfo_sCellInfo )";
            typeKind       = TECSTypeKind_DescriptorType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sCellInfo ))" );
            b_const        = false;
            b_volatile     = false;
            cSignatureInfo   = nTECSInfo_sCellInfoSignatureInfo.eSignatureInfo;
        };
        cell nTECSInfo::tPtrTypeInfo Descriptor_of_nTECSInfo_sRegionInfo_Ptr_TypeInfo{
            name           = "Descriptor( nTECSInfo_sRegionInfo )*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sRegionInfo )*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = Descriptor_of_nTECSInfo_sRegionInfoTypeInfo.eTypeInfo;
        };
        cell nTECSInfo::tDescriptorTypeInfo Descriptor_of_nTECSInfo_sRegionInfoTypeInfo{
            name           = "Descriptor( nTECSInfo_sRegionInfo )";
            typeKind       = TECSTypeKind_DescriptorType;
            size           = C_EXP( "sizeof(Descriptor( nTECSInfo_sRegionInfo ))" );
            b_const        = false;
            b_volatile     = false;
            cSignatureInfo   = nTECSInfo_sRegionInfoSignatureInfo.eSignatureInfo;
        };
        cell nTECSInfo::tPtrTypeInfo int_t_Ptr_TypeInfo{
            name           = "int_t*";
            typeKind       = TECSTypeKind_PtrType;
            size           = C_EXP( "sizeof(int_t*)" );
            b_const        = false;
            b_volatile     = false;
            cTypeInfo        = int_tTypeInfo.eTypeInfo;
        };

        /*** TECS information cell ***/
        cell nTECSInfo::tTECSInfoSub TECSInfoSub {
            cNamespaceInfo = _RootNamespaceInfo.eNamespaceInfo;
            cRegionInfo    = _LinkRootRegionInfo.eRegionInfo;
        } /* TECSInfoSub */;
    }; /* rTECSInfo */
};
