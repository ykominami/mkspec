import_C( "dupl-a.h" );  // dupl-b.h を include している
import_C( "dupl-b.h" );  // typedef int  INT;

typedef int32_t  INT32;
// typedef int32_t  INT32;
