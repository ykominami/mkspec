/*
 * simple なサンプル
 *
 * このサンプルは tecsgen/test/simple 階層に置いて実行する
 * Linux, Cygwin 環境で実行できるはず
 */
import_C( "cygwin_tecs.h" );

// ログ機能
import( <tSysLog.cdl> );
// カーネル機能
import( <cygwin_kernel.cdl> );
import( <rpc.cdl> );
import( <tSocketChannel.cdl> );
import( "tAlloc.cdl" );
import( "sSimple.cdl" );
import( "sSample.cdl" );

celltype tSimpleServer {
	require	tSysLog.eSysLog;
	entry	sSimple			eEnt;
/*	entry	sServerControl	eServerControl; */
};

[active]
celltype tSimpleClient {
	require	tSysLog.eSysLog;
	call	sSimple		cCall;
	/* call	sServerControl	cServerControl;	/* サーバをシャットダウンする */
	call	sSocketClientOpener	cOpener;	/* チャンネルを開く */
	call	sTask		cSampleTask;		/* */
	entry	sTaskBody	eMain;					/* メイン */
};


celltype tSampleServer {
	require	tSysLog.eSysLog;
	entry	sSample			eEnt;
};

[active]
celltype tSampleClient {
	require	tSysLog.eSysLog;
	call	sSample		cCall;
	/* call	sServerControl	cServerControl;	/* サーバをシャットダウンする */
	entry	sTaskBody	eMain;					/* メイン */
};

[out_through(),
 to_through(rServer ,SharedOpaqueRPCPlugin,
		"taskCelltype=tTask,PPAllocatorSize=1024,"
		"sharedChannelName= \"MyChannel\", "
		"substituteAllocator=\"Alloc.eAlloc=>CAlloc.eAlloc\", "   // 代替アロケータ指定
		"clientChannelCell= \"ClientChannel\", "
		"serverChannelCell= \"ServerChannel\" "
			), linkunit]
region rClient /*,nNamespace */ {
	cell tAlloc CAlloc {
	};
	cell tKernel KernelInClient {
	};
	cell tSysLog ClientSysLog {
	};
	cell tSocketClient ClientChannel {
	};
	[out_through(TracePlugin,"")]
//	[out_through()]
	region rCPon {
		cell tSimpleClient SimpleClient {
			cCall = rServer::rSPon::SimpleServer.eEnt;
			cSampleTask = Task1.eTask;
			cOpener = ClientChannel.eOpener;
		};
		cell tTask Task {
			cTaskBody = SimpleClient.eMain;
			priority = 1;
			stackSize = 4096;
			attribute = C_EXP( "TA_ACT" );
		};

	};
	cell tSampleClient SampleClient {
		cCall = rServer::SampleServer.eEnt;
	};
	cell tTask Task1 {
		cTaskBody = SampleClient.eMain;
		priority = 1;
		stackSize = 4096;
		attribute = C_EXP( "TA_NULL" );
	};
};

[in_through(), linkunit]
region rServer {
	cell	tSysLog	ServerSysLog {
	};
	cell tSocketServer ServerChannel {
	};

	// out_through() は TracePlugin から SysLog を参照するために必要
	[in_through(TracePlugin,""), out_through()]
//	[in_through(),out_through()]
	region rSPon {
		cell tAlloc Alloc {
		};
    //      cell tSysLog ServerSysLog {
    //      };
		cell tKernel KernelInServer {
		};
		[allocator(eEnt.func21.a=Alloc.eAlloc,
				   eEnt.func22.sta=Alloc.eAlloc,
				   eEnt.func23.str=Alloc.eAlloc,
				   eEnt.func24.msg=Alloc.eAlloc,
				   eEnt.func25.msg=Alloc.eAlloc,
				   eEnt.func26.sta=Alloc.eAlloc,
				   eEnt.func27.array2=Alloc.eAlloc,
				   eEnt.func31.a=Alloc.eAlloc,
				   eEnt.func32.sta=Alloc.eAlloc,
				   eEnt.func33.str=Alloc.eAlloc,
				   eEnt.func34.msg=Alloc.eAlloc,
				   eEnt.func35.msg=Alloc.eAlloc,
				   eEnt.func36.sta=Alloc.eAlloc,
				   eEnt.func37.sta=Alloc.eAlloc,
				   eEnt.func38.array2=Alloc.eAlloc,
				   eEnt.func39.arraySt=Alloc.eAlloc)]
		cell tSimpleServer SimpleServer {
		};
	};
	cell tSampleServer SampleServer { };
};

