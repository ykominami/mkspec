import( <cygwin_kernel.cdl> );
import( "HelloWorld.cdl" );
import( <TECSInfoAccessor.cdl> );

/*
 * TECSInfo 使用サンプル
 */
celltype tTaskMain {
    entry sTaskBody            eBody;
    call  nTECSInfo::sAccessor cAccessor;

    attr{
        int16_t NAME_LEN = 256;
    };
    var{
        [size_is(NAME_LEN)]
            char_t  *name;
        [size_is(NAME_LEN)]
            char_t  *name2;
    };
};


[in_through()]
region rTEMP{
    cell tTask Task {
        attribute = C_EXP("TA_ACT");
        priority      = 11;
        stackSize     = 4096;
        cTaskBody         = rTEMP::TaskMain.eBody;
    };
    cell tTaskMain TaskMain {
        cAccessor  = TECSInfoCompo.eAccessor;
    };

/******* TECSInfo cell *******/
    cell nTECSInfo::tTECSInfoCompo TECSInfoCompo {
        // cTECSInfo = rTECSInfo::TECSInfo.eTECSInfo;
        //  この結合は TECSInfoCompoPlugin により生成されるので結合不要
    };
};
