import_C( "cygwin_tecs.h" );
import( <cygwin_kernel.cdl> );
import( <utility.cdl> );

////// Signature Description //////
signature sHello {
	void  hello(void);
};

signature sTalkerSelector {
	void  getTalker([out]Descriptor(sHello) *talker, [in]int_t i);
	void  getNTalker([out]int_t *n);
};

////// Celltype Description //////
[singleton]
celltype tMainSingleArray {
	entry sTaskBody eMain;
	[ref_desc]
		call sHello cDefaultTalker;
	[dynamic]
		call sHello cTalker[];
	[dynamic,optional]
		call sHello cTalker2[2];
	call sTalkerSelector cTalkerSelector;
/*
    attr {
        int_t  a = 0;
    };
    var {
        int_t  v = 0;
    };
*/
};

[singleton]
celltype tMainSingleArrayForComp {
	entry sTaskBody eMain;
	[ref_desc]
		call sHello cDefaultTalker;
	[dynamic]
		call sHello cTalker[];
	[dynamic,optional]
		call sHello cTalker2[2];
	call sTalkerSelector cTalkerSelector;
/*
    attr {
        int_t  a = 0;
    };
    var {
        int_t  v = 0;
    };
*/
};

[singleton]
composite tCompMain {
	entry sTaskBody eMain;
	[ref_desc]
		call sHello cDefaultTalker;
	[dynamic]
		call sHello cTalker[];
	[dynamic,optional]
		call sHello cTalker2[2];
	call sTalkerSelector cTalkerSelector;
    cell tMainSingleArrayForComp Main {
        cDefaultTalker => composite.cDefaultTalker;
        cTalker => composite.cTalker;
        cTalker2 => composite.cTalker2;
        cTalkerSelector => composite.cTalkerSelector;
    };
    composite.eMain => Main.eMain;
};

celltype tTalkerSelector {
	entry sTalkerSelector eTalkerSelector;
	[ref_desc,optional]
		call  sHello  cHello[];
	attr {
		char_t *name = C_EXP( "\"$id$\"" );
	};
};

celltype tTalker {
	entry sHello eHello;
    attr {
        char_t *name = C_EXP( "\"$cell$\"" );
        char_t *message = "hello";
    };
};

////// Build Description //////
cell tSerialTask Task {
	cBodyArray[] = Main.eMain;
	cBodyArray[] = rComposite::CompMain.eMain;
	priority = 11;
	attribute = C_EXP( "TA_ACT" );
	stackSize = 256;
};

cell tMainSingleArray Main{
	cDefaultTalker = Talker0.eHello;
	cTalker[] = Talker0.eHello;
	cTalker[] = Talker1.eHello;
	cTalker[] = Talker2.eHello;
//	cTalker[] = Talker3.eHello;
	cTalkerSelector = Selector.eTalkerSelector;
};

cell tTalkerSelector Selector {
	cHello[0] = Talker0.eHello;
	cHello[1] = Talker1.eHello;
	cHello[2] = Talker2.eHello;
//	cHello[3] = Talker3.eHello;
	cHello[4] = Talker4.eHello;
	
};

cell tTalker Talker0 {};
cell tTalker Talker1 {};
cell tTalker Talker2 {};
//cell tTalker Talker3 {};
cell tTalker Talker4 {};

[in_through()]
region rComposite {
    cell tCompMain CompMain{
        cDefaultTalker = Talker0.eHello;
        cTalker[] = Talker0.eHello;
        cTalker[] = Talker1.eHello;
        cTalker[] = Talker2.eHello;
     //	cTalker[] = Talker3.eHello;
        cTalkerSelector = Selector.eTalkerSelector;
    };

    cell tTalkerSelector Selector {
        cHello[0] = Talker0.eHello;
        cHello[1] = Talker1.eHello;
        cHello[2] = Talker2.eHello;
     //	cHello[3] = Talker3.eHello;
        cHello[4] = Talker4.eHello;
    };

    cell tTalker Talker0 {};
    cell tTalker Talker1 {};
    cell tTalker Talker2 {};
//    cell tTalker Talker3 {};
    cell tTalker Talker4 {};
};


