import( "cygwin_kernel.cdl" );
import( "tSysLog.cdl" );
cell tSysLog SysLog {};
cell tKernel Kernel {};

[deviate]
signature sAlloc {
  ER  alloc( [in]int32_t size, [out]void **p );
  ER  dealloc( [in]const void *p );
};
celltype tAlloc {
  entry sAlloc eA;
  attr {
    int32_t  size = 8192;
  };
  var {
    [size_is(size)]
    int8_t  *buffer;
  };
};

cell tAlloc alloc {
};

signature sSendRecv {
  /* この関数名に send, receive を使ってしまうと allocator 指定できない */
  ER snd( [send(sAlloc),size_is(sz)]int8_t *buf, [in]int32_t  sz );
  ER rcv( [receive(sAlloc),size_is(*sz)]int8_t **buf, [out]int32_t  *sz );
};

/****  Server Celltypes ****/
celltype tTestComponent {
  entry  sSendRecv eS;
  entry  sSendRecv eA[2];
};

celltype tTestComponent2 {
  entry  sSendRecv eS;
  entry  sSendRecv eA[];
};

composite tTestComponent3{
  entry  sSendRecv eS;
  entry  sSendRecv eA[];

  cell tTestComponent2 Cell {
  };
  composite.eS => Cell.eS;
  composite.eA => Cell.eA;
};

/****  Server Cells ****/
[allocator(
   eS.snd.buf=alloc.eA,
   eS.rcv.buf=alloc.eA,
   eA[0].snd.buf=alloc.eA,
   eA[1].snd.buf=alloc.eA,
   eA[0].rcv.buf=alloc.eA,
   eA[1].rcv.buf=alloc.eA
)]
cell tTestComponent Comp{
};

[allocator(
   eS.snd.buf=alloc.eA,
   eS.rcv.buf=alloc.eA,
   eA[0].snd.buf=alloc.eA,
   eA[1].snd.buf=alloc.eA,
   eA[0].rcv.buf=alloc.eA,
   eA[1].rcv.buf=alloc.eA
)]
cell tTestComponent3 Comp2{
};

/**** Client Celltype ****/
celltype tTestClient {
    [omit]
        call   sSendRecv cS;
    [omit]
        call   sSendRecv cA[2];
    entry  sTaskBody eBody;
};

cell tTestClient Cl {
  cS    = Comp.eS;
  cA[0] = Comp.eA[0];
  cA[1] = Comp.eA[1];
};


composite tTestClient2 {
    [omit]
        call   sSendRecv cS;
    [omit]
        call   sSendRecv cA[2];
    entry  sTaskBody eBody;
    cell tTestClient Cell {
        cS    => composite.cS;
        cA    => composite.cA;
    };
    composite.eBody => Cell.eBody;
    
};

cell tTestClient2 Cl2 {
  [through(TracePlugin,"")]
  cS =    Comp2.eS;
  cA[0] = Comp2.eA[0];
  cA[1] = Comp2.eA[1];
};

cell tTask Task1{
    attribute = C_EXP("TA_ACT");
    priority = 15;
	stackSize = 4096;
    cTaskBody = Cl.eBody;
};

cell tTask Task2{
    attribute = C_EXP("TA_ACT");
    priority = 15;
	stackSize = 4096;
    cTaskBody = Cl2.eBody;
};
