import_C( "cygwin_syslog.h" );
