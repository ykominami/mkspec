signature sSample {
	void	func(void);
};
